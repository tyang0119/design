
module pipe ( clk, reset, A, B, result, wrAddr );
  input [15:0] A;
  input [15:0] B;
  output [15:0] result;
  input [3:0] wrAddr;
  input clk, reset;
  wire   \nextState[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n528, n529, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n602, n603, n604, n605,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232;
  wire   [8:0] aAQ;
  wire   [15:0] doA;
  wire   [8:0] aBQ;
  wire   [15:0] doB;
  wire   [15:0] ramAQ;
  wire   [15:0] ramBQ;
  wire   [15:0] result2;
  wire   [15:0] partialQ;
  wire   [15:0] multQ;
  wire   [15:0] counterQ;
  wire   [1:0] state;
  wire   [3:0] \mult/state ;
  wire   [6:0] \mult/counterQ ;
  wire   [31:0] \mult/productQ ;
  wire   [31:0] \mult/storeQ ;

  ramA_2 ramA ( .clk(clk), .we(\nextState[0] ), .a(aAQ), .di(A), .do(doA) );
  ramB_2 ramB ( .clk(clk), .we(\nextState[0] ), .a(aBQ), .di(B), .do(doB) );
  dp_1 \state_reg[0]  ( .ip(n684), .ck(clk), .q(state[0]) );
  dp_1 \state_reg[1]  ( .ip(n683), .ck(clk), .q(state[1]) );
  dp_1 \ramAQ_reg[15]  ( .ip(n682), .ck(clk), .q(ramAQ[15]) );
  dp_1 \ramAQ_reg[13]  ( .ip(n680), .ck(clk), .q(ramAQ[13]) );
  dp_1 \ramAQ_reg[12]  ( .ip(n679), .ck(clk), .q(ramAQ[12]) );
  dp_1 \ramAQ_reg[11]  ( .ip(n678), .ck(clk), .q(ramAQ[11]) );
  dp_1 \ramAQ_reg[10]  ( .ip(n677), .ck(clk), .q(ramAQ[10]) );
  dp_1 \ramAQ_reg[7]  ( .ip(n674), .ck(clk), .q(ramAQ[7]) );
  dp_1 \ramAQ_reg[6]  ( .ip(n673), .ck(clk), .q(ramAQ[6]) );
  dp_1 \ramAQ_reg[5]  ( .ip(n672), .ck(clk), .q(ramAQ[5]) );
  dp_1 \ramAQ_reg[0]  ( .ip(n667), .ck(clk), .q(ramAQ[0]) );
  dp_1 \ramBQ_reg[15]  ( .ip(n666), .ck(clk), .q(ramBQ[15]) );
  dp_1 \ramBQ_reg[14]  ( .ip(n665), .ck(clk), .q(ramBQ[14]) );
  dp_1 \ramBQ_reg[13]  ( .ip(n664), .ck(clk), .q(ramBQ[13]) );
  dp_1 \ramBQ_reg[12]  ( .ip(n663), .ck(clk), .q(ramBQ[12]) );
  dp_1 \ramBQ_reg[11]  ( .ip(n662), .ck(clk), .q(ramBQ[11]) );
  dp_1 \ramBQ_reg[10]  ( .ip(n661), .ck(clk), .q(ramBQ[10]) );
  dp_1 \ramBQ_reg[9]  ( .ip(n660), .ck(clk), .q(ramBQ[9]) );
  dp_1 \ramBQ_reg[8]  ( .ip(n659), .ck(clk), .q(ramBQ[8]) );
  dp_1 \ramBQ_reg[6]  ( .ip(n657), .ck(clk), .q(ramBQ[6]) );
  dp_1 \ramBQ_reg[5]  ( .ip(n656), .ck(clk), .q(ramBQ[5]) );
  dp_1 \ramBQ_reg[4]  ( .ip(n655), .ck(clk), .q(ramBQ[4]) );
  dp_1 \ramBQ_reg[3]  ( .ip(n654), .ck(clk), .q(ramBQ[3]) );
  dp_1 \ramBQ_reg[2]  ( .ip(n653), .ck(clk), .q(ramBQ[2]) );
  dp_1 \ramBQ_reg[1]  ( .ip(n652), .ck(clk), .q(ramBQ[1]) );
  dp_1 \ramBQ_reg[0]  ( .ip(n651), .ck(clk), .q(ramBQ[0]) );
  dp_1 \counterQ_reg[0]  ( .ip(n650), .ck(clk), .q(counterQ[0]) );
  dp_1 \partialQ_reg[1]  ( .ip(n544), .ck(clk), .q(partialQ[1]) );
  dp_1 \partialQ_reg[2]  ( .ip(n543), .ck(clk), .q(partialQ[2]) );
  dp_1 \partialQ_reg[3]  ( .ip(n542), .ck(clk), .q(partialQ[3]) );
  dp_1 \partialQ_reg[4]  ( .ip(n541), .ck(clk), .q(partialQ[4]) );
  dp_1 \partialQ_reg[5]  ( .ip(n540), .ck(clk), .q(partialQ[5]) );
  dp_1 \partialQ_reg[6]  ( .ip(n539), .ck(clk), .q(partialQ[6]) );
  dp_1 \partialQ_reg[7]  ( .ip(n538), .ck(clk), .q(partialQ[7]) );
  dp_1 \partialQ_reg[9]  ( .ip(n536), .ck(clk), .q(partialQ[9]) );
  dp_1 \partialQ_reg[12]  ( .ip(n533), .ck(clk), .q(partialQ[12]) );
  dp_1 \mult/state_reg[1]  ( .ip(n634), .ck(clk), .q(\mult/state [1]) );
  dp_1 \mult/storeQ_reg[17]  ( .ip(n2231), .ck(clk), .q(\mult/storeQ [17]) );
  dp_1 \mult/storeQ_reg[21]  ( .ip(n604), .ck(clk), .q(\mult/storeQ [21]) );
  dp_1 \mult/storeQ_reg[7]  ( .ip(n618), .ck(clk), .q(\mult/storeQ [7]) );
  dp_1 \mult/storeQ_reg[23]  ( .ip(n602), .ck(clk), .q(\mult/storeQ [23]) );
  dp_1 \mult/storeQ_reg[15]  ( .ip(n610), .ck(clk), .q(\mult/storeQ [15]) );
  dp_1 \mult/storeQ_reg[19]  ( .ip(n2230), .ck(clk), .q(\mult/storeQ [19]) );
  dp_1 \mult/storeQ_reg[6]  ( .ip(n619), .ck(clk), .q(\mult/storeQ [6]) );
  dp_1 \mult/storeQ_reg[22]  ( .ip(n603), .ck(clk), .q(\mult/storeQ [22]) );
  dp_1 \mult/storeQ_reg[18]  ( .ip(n2229), .ck(clk), .q(\mult/storeQ [18]) );
  dp_1 \mult/storeQ_reg[4]  ( .ip(n621), .ck(clk), .q(\mult/storeQ [4]) );
  dp_1 \mult/storeQ_reg[20]  ( .ip(n605), .ck(clk), .q(\mult/storeQ [20]) );
  dp_1 \mult/storeQ_reg[8]  ( .ip(n617), .ck(clk), .q(\mult/storeQ [8]) );
  dp_1 \mult/storeQ_reg[16]  ( .ip(n609), .ck(clk), .q(\mult/storeQ [16]) );
  dp_1 \mult/storeQ_reg[0]  ( .ip(n625), .ck(clk), .q(\mult/storeQ [0]) );
  dp_1 \mult/productQ_reg[0]  ( .ip(n593), .ck(clk), .q(\mult/productQ [0]) );
  dp_1 \mult/productQ_reg[4]  ( .ip(n589), .ck(clk), .q(\mult/productQ [4]) );
  dp_1 \mult/productQ_reg[7]  ( .ip(n586), .ck(clk), .q(\mult/productQ [7]) );
  dp_1 \mult/productQ_reg[20]  ( .ip(n573), .ck(clk), .q(\mult/productQ [20])
         );
  dp_1 \mult/productQ_reg[22]  ( .ip(n571), .ck(clk), .q(\mult/productQ [22])
         );
  dp_1 \multQ_reg[0]  ( .ip(n561), .ck(clk), .q(multQ[0]) );
  dp_1 \multQ_reg[1]  ( .ip(n560), .ck(clk), .q(multQ[1]) );
  dp_1 \multQ_reg[2]  ( .ip(n559), .ck(clk), .q(multQ[2]) );
  dp_1 \multQ_reg[3]  ( .ip(n558), .ck(clk), .q(multQ[3]) );
  dp_1 \multQ_reg[5]  ( .ip(n556), .ck(clk), .q(multQ[5]) );
  dp_1 \multQ_reg[6]  ( .ip(n555), .ck(clk), .q(multQ[6]) );
  dp_1 \multQ_reg[7]  ( .ip(n554), .ck(clk), .q(multQ[7]) );
  dp_1 \multQ_reg[8]  ( .ip(n553), .ck(clk), .q(multQ[8]) );
  dp_1 \multQ_reg[9]  ( .ip(n552), .ck(clk), .q(multQ[9]) );
  dp_1 \multQ_reg[10]  ( .ip(n551), .ck(clk), .q(multQ[10]) );
  dp_1 \multQ_reg[11]  ( .ip(n550), .ck(clk), .q(multQ[11]) );
  dp_1 \multQ_reg[12]  ( .ip(n549), .ck(clk), .q(multQ[12]) );
  dp_1 \multQ_reg[14]  ( .ip(n547), .ck(clk), .q(multQ[14]) );
  dp_1 \multQ_reg[15]  ( .ip(n546), .ck(clk), .q(multQ[15]) );
  dp_1 \aBQ_reg[0]  ( .ip(n18), .ck(clk), .q(aBQ[0]) );
  dp_1 \aBQ_reg[8]  ( .ip(n17), .ck(clk), .q(aBQ[8]) );
  dp_1 \aAQ_reg[8]  ( .ip(n16), .ck(clk), .q(aAQ[8]) );
  dp_1 \aAQ_reg[7]  ( .ip(n15), .ck(clk), .q(aAQ[7]) );
  dp_1 \aAQ_reg[6]  ( .ip(n14), .ck(clk), .q(aAQ[6]) );
  dp_1 \aAQ_reg[5]  ( .ip(n13), .ck(clk), .q(aAQ[5]) );
  dp_1 \aAQ_reg[4]  ( .ip(n12), .ck(clk), .q(aAQ[4]) );
  dp_1 \aAQ_reg[3]  ( .ip(n11), .ck(clk), .q(aAQ[3]) );
  dp_1 \aAQ_reg[2]  ( .ip(n10), .ck(clk), .q(aAQ[2]) );
  dp_1 \aAQ_reg[1]  ( .ip(n9), .ck(clk), .q(aAQ[1]) );
  dp_1 \aAQ_reg[0]  ( .ip(n8), .ck(clk), .q(aAQ[0]) );
  dp_1 \aBQ_reg[7]  ( .ip(n7), .ck(clk), .q(aBQ[7]) );
  dp_1 \aBQ_reg[6]  ( .ip(n6), .ck(clk), .q(aBQ[6]) );
  dp_1 \aBQ_reg[5]  ( .ip(n5), .ck(clk), .q(aBQ[5]) );
  dp_1 \aBQ_reg[4]  ( .ip(n4), .ck(clk), .q(aBQ[4]) );
  dp_1 \aBQ_reg[3]  ( .ip(n3), .ck(clk), .q(aBQ[3]) );
  dp_1 \aBQ_reg[2]  ( .ip(n2), .ck(clk), .q(aBQ[2]) );
  dp_2 \counterQ_reg[2]  ( .ip(n648), .ck(clk), .q(counterQ[2]) );
  dp_2 \counterQ_reg[6]  ( .ip(n644), .ck(clk), .q(counterQ[6]) );
  dp_2 \counterQ_reg[10]  ( .ip(n640), .ck(clk), .q(counterQ[10]) );
  dp_2 \counterQ_reg[12]  ( .ip(n638), .ck(clk), .q(counterQ[12]) );
  dp_2 \counterQ_reg[1]  ( .ip(n649), .ck(clk), .q(counterQ[1]) );
  dp_2 \counterQ_reg[4]  ( .ip(n646), .ck(clk), .q(counterQ[4]) );
  dp_2 \counterQ_reg[8]  ( .ip(n642), .ck(clk), .q(counterQ[8]) );
  nand2_1 U710 ( .ip1(n528), .ip2(n529), .op(\nextState[0] ) );
  dp_4 \mult/counterQ_reg[2]  ( .ip(n628), .ck(clk), .q(\mult/counterQ [2]) );
  dp_2 \mult/productQ_reg[12]  ( .ip(n581), .ck(clk), .q(\mult/productQ [12])
         );
  dp_2 \mult/storeQ_reg[12]  ( .ip(n613), .ck(clk), .q(\mult/storeQ [12]) );
  lp_1 \mult/PRODUCT_reg[5]  ( .ck(n1273), .ip(\mult/productQ [13]), .q(
        result2[5]) );
  dp_2 \mult/productQ_reg[3]  ( .ip(n590), .ck(clk), .q(\mult/productQ [3]) );
  lp_1 \mult/PRODUCT_reg[2]  ( .ck(n1273), .ip(\mult/productQ [10]), .q(
        result2[2]) );
  lp_1 \mult/PRODUCT_reg[1]  ( .ck(n1273), .ip(\mult/productQ [9]), .q(
        result2[1]) );
  dp_2 \mult/productQ_reg[14]  ( .ip(n579), .ck(clk), .q(\mult/productQ [14])
         );
  dp_2 \mult/storeQ_reg[14]  ( .ip(n611), .ck(clk), .q(\mult/storeQ [14]) );
  lp_1 \mult/PRODUCT_reg[4]  ( .ck(n1273), .ip(\mult/productQ [12]), .q(
        result2[4]) );
  dp_2 \mult/storeQ_reg[11]  ( .ip(n614), .ck(clk), .q(\mult/storeQ [11]) );
  dp_2 \mult/productQ_reg[11]  ( .ip(n582), .ck(clk), .q(\mult/productQ [11])
         );
  dp_2 \mult/state_reg[0]  ( .ip(n632), .ck(clk), .q(\mult/state [0]) );
  dp_2 \mult/counterQ_reg[0]  ( .ip(n626), .ck(clk), .q(\mult/counterQ [0]) );
  dp_2 \mult/productQ_reg[13]  ( .ip(n580), .ck(clk), .q(\mult/productQ [13])
         );
  dp_2 \mult/counterQ_reg[1]  ( .ip(n627), .ck(clk), .q(\mult/counterQ [1]) );
  dp_2 \mult/storeQ_reg[13]  ( .ip(n612), .ck(clk), .q(\mult/storeQ [13]) );
  lp_1 \mult/PRODUCT_reg[13]  ( .ck(n1273), .ip(\mult/productQ [21]), .q(
        result2[13]) );
  dp_2 \mult/storeQ_reg[3]  ( .ip(n622), .ck(clk), .q(\mult/storeQ [3]) );
  dp_2 \counterQ_reg[9]  ( .ip(n641), .ck(clk), .q(counterQ[9]) );
  dp_2 \mult/productQ_reg[2]  ( .ip(n591), .ck(clk), .q(\mult/productQ [2]) );
  dp_2 \mult/storeQ_reg[2]  ( .ip(n623), .ck(clk), .q(\mult/storeQ [2]) );
  dp_2 \mult/storeQ_reg[1]  ( .ip(n624), .ck(clk), .q(\mult/storeQ [1]) );
  dp_2 \mult/productQ_reg[10]  ( .ip(n583), .ck(clk), .q(\mult/productQ [10])
         );
  dp_2 \mult/productQ_reg[15]  ( .ip(n578), .ck(clk), .q(\mult/productQ [15])
         );
  dp_2 \mult/productQ_reg[1]  ( .ip(n592), .ck(clk), .q(\mult/productQ [1]) );
  dp_2 \mult/counterQ_reg[3]  ( .ip(n629), .ck(clk), .q(\mult/counterQ [3]) );
  dp_2 \mult/productQ_reg[8]  ( .ip(n585), .ck(clk), .q(\mult/productQ [8]) );
  dp_2 \mult/storeQ_reg[9]  ( .ip(n616), .ck(clk), .q(\mult/storeQ [9]) );
  dp_2 \counterQ_reg[11]  ( .ip(n639), .ck(clk), .q(counterQ[11]) );
  dp_2 \ramAQ_reg[8]  ( .ip(n675), .ck(clk), .q(ramAQ[8]) );
  dp_2 \ramAQ_reg[2]  ( .ip(n669), .ck(clk), .q(ramAQ[2]) );
  lp_1 \result_reg[13]  ( .ck(n2232), .ip(partialQ[13]), .q(result[13]) );
  lp_1 \result_reg[8]  ( .ck(n2232), .ip(partialQ[8]), .q(result[8]) );
  lp_1 \result_reg[5]  ( .ck(n2232), .ip(partialQ[5]), .q(result[5]) );
  lp_1 \result_reg[10]  ( .ck(n2232), .ip(partialQ[10]), .q(result[10]) );
  lp_1 \result_reg[7]  ( .ck(n2232), .ip(partialQ[7]), .q(result[7]) );
  lp_1 \result_reg[9]  ( .ck(n2232), .ip(partialQ[9]), .q(result[9]) );
  lp_1 \result_reg[1]  ( .ck(n2232), .ip(partialQ[1]), .q(result[1]) );
  lp_1 \result_reg[2]  ( .ck(n2232), .ip(partialQ[2]), .q(result[2]) );
  lp_1 \result_reg[3]  ( .ck(n2232), .ip(partialQ[3]), .q(result[3]) );
  lp_1 \result_reg[4]  ( .ck(n2232), .ip(partialQ[4]), .q(result[4]) );
  lp_1 \result_reg[11]  ( .ck(n2232), .ip(partialQ[11]), .q(result[11]) );
  lp_1 \result_reg[12]  ( .ck(n2232), .ip(partialQ[12]), .q(result[12]) );
  lp_1 \result_reg[14]  ( .ck(n2232), .ip(partialQ[14]), .q(result[14]) );
  lp_1 \result_reg[15]  ( .ck(n2232), .ip(partialQ[15]), .q(result[15]) );
  lp_1 \result_reg[6]  ( .ck(n2232), .ip(partialQ[6]), .q(result[6]) );
  lp_1 \result_reg[0]  ( .ck(n2232), .ip(partialQ[0]), .q(result[0]) );
  lp_1 \mult/PRODUCT_reg[7]  ( .ck(n1273), .ip(\mult/productQ [15]), .q(
        result2[7]) );
  lp_1 \mult/PRODUCT_reg[15]  ( .ck(n1273), .ip(\mult/productQ [23]), .q(
        result2[15]) );
  lp_1 \mult/PRODUCT_reg[0]  ( .ck(n1273), .ip(\mult/productQ [8]), .q(
        result2[0]) );
  lp_1 \mult/PRODUCT_reg[3]  ( .ck(n1273), .ip(\mult/productQ [11]), .q(
        result2[3]) );
  lp_1 \mult/PRODUCT_reg[6]  ( .ck(n1273), .ip(\mult/productQ [14]), .q(
        result2[6]) );
  lp_1 \mult/PRODUCT_reg[14]  ( .ck(n1273), .ip(\mult/productQ [22]), .q(
        result2[14]) );
  lp_1 \mult/PRODUCT_reg[8]  ( .ck(n1273), .ip(\mult/productQ [16]), .q(
        result2[8]) );
  lp_1 \mult/PRODUCT_reg[9]  ( .ck(n1273), .ip(\mult/productQ [17]), .q(
        result2[9]) );
  lp_1 \mult/PRODUCT_reg[10]  ( .ck(n1273), .ip(\mult/productQ [18]), .q(
        result2[10]) );
  lp_1 \mult/PRODUCT_reg[11]  ( .ck(n1273), .ip(\mult/productQ [19]), .q(
        result2[11]) );
  lp_1 \mult/PRODUCT_reg[12]  ( .ck(n1273), .ip(\mult/productQ [20]), .q(
        result2[12]) );
  dp_2 \mult/counterQ_reg[4]  ( .ip(n630), .ck(clk), .q(\mult/counterQ [4]) );
  dp_2 \mult/productQ_reg[9]  ( .ip(n584), .ck(clk), .q(\mult/productQ [9]) );
  dp_2 \partialQ_reg[11]  ( .ip(n534), .ck(clk), .q(partialQ[11]) );
  dp_2 \multQ_reg[4]  ( .ip(n557), .ck(clk), .q(multQ[4]) );
  dksp_1 \partialQ_reg[15]  ( .ip(n2159), .sb(n2160), .ck(clk), .q(
        partialQ[15]), .qb() );
  dp_2 \partialQ_reg[13]  ( .ip(n532), .ck(clk), .q(partialQ[13]) );
  dp_2 \mult/storeQ_reg[10]  ( .ip(n615), .ck(clk), .q(\mult/storeQ [10]) );
  dp_2 \counterQ_reg[5]  ( .ip(n645), .ck(clk), .q(counterQ[5]) );
  dp_2 \mult/productQ_reg[5]  ( .ip(n588), .ck(clk), .q(\mult/productQ [5]) );
  dp_2 \mult/storeQ_reg[5]  ( .ip(n620), .ck(clk), .q(\mult/storeQ [5]) );
  dp_2 \counterQ_reg[14]  ( .ip(n636), .ck(clk), .q(counterQ[14]) );
  dp_2 \counterQ_reg[15]  ( .ip(n635), .ck(clk), .q(counterQ[15]) );
  dp_2 \partialQ_reg[10]  ( .ip(n535), .ck(clk), .q(partialQ[10]) );
  dp_2 \counterQ_reg[13]  ( .ip(n637), .ck(clk), .q(counterQ[13]) );
  dp_2 \partialQ_reg[14]  ( .ip(n531), .ck(clk), .q(partialQ[14]) );
  dp_2 \partialQ_reg[0]  ( .ip(n545), .ck(clk), .q(partialQ[0]) );
  dp_2 \partialQ_reg[8]  ( .ip(n537), .ck(clk), .q(partialQ[8]) );
  dp_2 \counterQ_reg[7]  ( .ip(n643), .ck(clk), .q(counterQ[7]) );
  dp_2 \aBQ_reg[1]  ( .ip(n1), .ck(clk), .q(aBQ[1]) );
  drp_1 \counterQ_reg[3]  ( .ip(n647), .ck(clk), .rb(1'b1), .q(counterQ[3]) );
  dp_2 \mult/counterQ_reg[5]  ( .ip(n631), .ck(clk), .q(\mult/counterQ [5]) );
  dp_1 \ramAQ_reg[1]  ( .ip(n668), .ck(clk), .q(ramAQ[1]) );
  dp_1 \ramBQ_reg[7]  ( .ip(n658), .ck(clk), .q(ramBQ[7]) );
  dp_2 \mult/productQ_reg[21]  ( .ip(n572), .ck(clk), .q(\mult/productQ [21])
         );
  dp_2 \mult/productQ_reg[6]  ( .ip(n587), .ck(clk), .q(\mult/productQ [6]) );
  dp_2 \mult/productQ_reg[16]  ( .ip(n577), .ck(clk), .q(\mult/productQ [16])
         );
  dp_2 \mult/productQ_reg[19]  ( .ip(n574), .ck(clk), .q(\mult/productQ [19])
         );
  dp_2 \mult/productQ_reg[17]  ( .ip(n576), .ck(clk), .q(\mult/productQ [17])
         );
  dp_2 \mult/productQ_reg[18]  ( .ip(n575), .ck(clk), .q(\mult/productQ [18])
         );
  dp_2 \mult/productQ_reg[23]  ( .ip(n570), .ck(clk), .q(\mult/productQ [23])
         );
  dp_1 \ramAQ_reg[3]  ( .ip(n670), .ck(clk), .q(ramAQ[3]) );
  dp_1 \multQ_reg[13]  ( .ip(n548), .ck(clk), .q(multQ[13]) );
  dp_1 \ramAQ_reg[14]  ( .ip(n681), .ck(clk), .q(ramAQ[14]) );
  dp_1 \ramAQ_reg[9]  ( .ip(n676), .ck(clk), .q(ramAQ[9]) );
  dp_1 \ramAQ_reg[4]  ( .ip(n671), .ck(clk), .q(ramAQ[4]) );
  buf_2 U711 ( .ip(n1856), .op(n2151) );
  inv_2 U712 ( .ip(n1795), .op(n2092) );
  inv_2 U713 ( .ip(n1736), .op(n721) );
  buf_2 U714 ( .ip(n1354), .op(n2059) );
  inv_2 U715 ( .ip(n1219), .op(n1201) );
  inv_4 U716 ( .ip(n1917), .op(n1293) );
  buf_2 U717 ( .ip(n805), .op(n2069) );
  buf_2 U718 ( .ip(n1354), .op(n2049) );
  inv_2 U719 ( .ip(n805), .op(n1354) );
  inv_2 U720 ( .ip(n1976), .op(n2081) );
  nand2_2 U721 ( .ip1(n1150), .ip2(partialQ[12]), .op(n2016) );
  inv_2 U722 ( .ip(\mult/counterQ [3]), .op(n1976) );
  nand2_2 U723 ( .ip1(n694), .ip2(n693), .op(n696) );
  nor2_2 U724 ( .ip1(n1470), .ip2(n1469), .op(n1471) );
  inv_4 U725 ( .ip(n1727), .op(n1736) );
  and2_2 U726 ( .ip1(n873), .ip2(n872), .op(n2074) );
  nor2_2 U727 ( .ip1(n868), .ip2(n867), .op(n873) );
  inv_2 U728 ( .ip(n2077), .op(n2078) );
  inv_2 U729 ( .ip(n1727), .op(n2077) );
  inv_2 U730 ( .ip(n1736), .op(n1805) );
  nand2_4 U731 ( .ip1(n1220), .ip2(n1201), .op(n1795) );
  nor3_2 U732 ( .ip1(n1779), .ip2(n1778), .ip3(n1777), .op(n1780) );
  nand2_2 U733 ( .ip1(n1776), .ip2(n1775), .op(n1777) );
  nor2_2 U734 ( .ip1(n2069), .ip2(n1888), .op(n1881) );
  inv_2 U735 ( .ip(partialQ[3]), .op(n787) );
  inv_2 U736 ( .ip(n1132), .op(n1872) );
  nand2_2 U737 ( .ip1(n1135), .ip2(partialQ[11]), .op(n1873) );
  inv_2 U738 ( .ip(partialQ[10]), .op(n1918) );
  inv_1 U739 ( .ip(n689), .op(n1922) );
  nand2_1 U740 ( .ip1(n1918), .ip2(n1239), .op(n689) );
  nand3_2 U741 ( .ip1(n1709), .ip2(n799), .ip3(n1699), .op(n2013) );
  nand2_2 U742 ( .ip1(n1239), .ip2(n1918), .op(n1144) );
  nand2_2 U743 ( .ip1(n1145), .ip2(n1144), .op(n1876) );
  nand2_1 U744 ( .ip1(n1232), .ip2(n1231), .op(n1233) );
  nand2_2 U745 ( .ip1(n773), .ip2(n787), .op(n772) );
  nand2_2 U746 ( .ip1(n1481), .ip2(n772), .op(n1501) );
  nand2_1 U747 ( .ip1(n1226), .ip2(n1227), .op(n1504) );
  nand2_1 U748 ( .ip1(n1749), .ip2(n1745), .op(n1227) );
  inv_2 U749 ( .ip(n1233), .op(n1499) );
  nand2_2 U750 ( .ip1(n1234), .ip2(n1499), .op(n1865) );
  nand2_2 U751 ( .ip1(n788), .ip2(n787), .op(n1231) );
  nand2_1 U752 ( .ip1(n690), .ip2(n765), .op(n763) );
  nor2_1 U753 ( .ip1(n761), .ip2(n760), .op(n690) );
  nor2_2 U754 ( .ip1(n691), .ip2(n895), .op(n897) );
  nor2_2 U755 ( .ip1(n932), .ip2(n893), .op(n691) );
  nand2_1 U756 ( .ip1(n753), .ip2(n692), .op(n756) );
  nor2_2 U757 ( .ip1(counterQ[6]), .ip2(counterQ[2]), .op(n692) );
  inv_4 U758 ( .ip(n696), .op(n1618) );
  inv_1 U759 ( .ip(\mult/counterQ [1]), .op(n693) );
  inv_1 U760 ( .ip(\mult/counterQ [0]), .op(n694) );
  nor2_1 U761 ( .ip1(n1649), .ip2(n998), .op(n1811) );
  nand2_1 U762 ( .ip1(aBQ[3]), .ip2(aBQ[2]), .op(n2196) );
  inv_1 U763 ( .ip(partialQ[8]), .op(n1700) );
  inv_1 U764 ( .ip(n1785), .op(n1978) );
  nand2_1 U765 ( .ip1(n1208), .ip2(n1354), .op(n1216) );
  or3_1 U766 ( .ip1(n1786), .ip2(n1802), .ip3(n1575), .op(n695) );
  or2_1 U767 ( .ip1(n2062), .ip2(n2061), .op(n697) );
  nand2_1 U768 ( .ip1(n764), .ip2(n1227), .op(n770) );
  nand2_1 U769 ( .ip1(n698), .ip2(n1160), .op(n1161) );
  inv_1 U770 ( .ip(n1211), .op(n698) );
  nand2_1 U771 ( .ip1(n1158), .ip2(n699), .op(n1211) );
  inv_1 U772 ( .ip(n700), .op(n699) );
  nand2_1 U773 ( .ip1(n2022), .ip2(n1157), .op(n700) );
  nand2_1 U774 ( .ip1(n1354), .ip2(n1710), .op(n1705) );
  nand2_1 U775 ( .ip1(n1701), .ip2(n1702), .op(n1710) );
  nand2_1 U776 ( .ip1(n1613), .ip2(ramBQ[6]), .op(n823) );
  nand2_1 U777 ( .ip1(n1228), .ip2(n1466), .op(n1498) );
  nand2_1 U778 ( .ip1(n795), .ip2(n1266), .op(n1228) );
  nand2_1 U779 ( .ip1(n1573), .ip2(n701), .op(n605) );
  nand2_1 U780 ( .ip1(n1571), .ip2(n1572), .op(n701) );
  nand3_1 U781 ( .ip1(n815), .ip2(n816), .ip3(n811), .op(n536) );
  nand2_1 U782 ( .ip1(n702), .ip2(n917), .op(n920) );
  inv_1 U783 ( .ip(n703), .op(n702) );
  nand2_1 U784 ( .ip1(n915), .ip2(n719), .op(n703) );
  nand2_1 U785 ( .ip1(n1906), .ip2(n704), .op(n1913) );
  nand3_1 U786 ( .ip1(n1902), .ip2(n1903), .ip3(n1904), .op(n704) );
  nand2_1 U787 ( .ip1(n707), .ip2(n705), .op(n1564) );
  inv_1 U788 ( .ip(n706), .op(n705) );
  nand2_1 U789 ( .ip1(n1976), .ip2(n1793), .op(n706) );
  inv_1 U790 ( .ip(n1730), .op(n707) );
  buf_4 U791 ( .ip(n1624), .op(n708) );
  nand3_1 U792 ( .ip1(n697), .ip2(n2072), .ip3(n709), .op(n539) );
  nor2_1 U793 ( .ip1(n710), .ip2(n2063), .op(n709) );
  inv_1 U794 ( .ip(n711), .op(n710) );
  nand2_1 U795 ( .ip1(partialQ[6]), .ip2(n2064), .op(n711) );
  nor2_2 U796 ( .ip1(n2016), .ip2(n1152), .op(n1153) );
  or3_2 U797 ( .ip1(n798), .ip2(n797), .ip3(n796), .op(n1709) );
  nand2_1 U798 ( .ip1(\mult/storeQ [15]), .ip2(n1727), .op(n722) );
  nand2_2 U799 ( .ip1(n876), .ip2(n1529), .op(n1220) );
  inv_1 U800 ( .ip(n1746), .op(n713) );
  xor2_2 U801 ( .ip1(n2006), .ip2(n1400), .op(n737) );
  nor2_1 U802 ( .ip1(n2161), .ip2(n2216), .op(n2221) );
  nor2_1 U803 ( .ip1(n2161), .ip2(n2200), .op(n2205) );
  nor3_1 U804 ( .ip1(n1082), .ip2(n1081), .ip3(n1080), .op(n1083) );
  nor2_1 U805 ( .ip1(n1408), .ip2(n1423), .op(n1417) );
  inv_4 U806 ( .ip(n1311), .op(n1387) );
  nor2_1 U807 ( .ip1(n2115), .ip2(n1825), .op(n2145) );
  nand2_2 U808 ( .ip1(aAQ[3]), .ip2(aAQ[2]), .op(n2212) );
  nand2_1 U809 ( .ip1(n723), .ip2(n722), .op(n610) );
  nand2_1 U810 ( .ip1(n1271), .ip2(n1270), .op(n544) );
  xnor2_1 U811 ( .ip1(n1490), .ip2(n1489), .op(n1491) );
  and2_1 U812 ( .ip1(n810), .ip2(n809), .op(n811) );
  nand2_1 U813 ( .ip1(n726), .ip2(n725), .op(n724) );
  nand2_1 U814 ( .ip1(n1791), .ip2(n1790), .op(n725) );
  nor3_1 U815 ( .ip1(n1978), .ip2(n1673), .ip3(n1672), .op(n1674) );
  nor2_1 U816 ( .ip1(n2132), .ip2(n2131), .op(n2133) );
  nor3_1 U817 ( .ip1(n1693), .ip2(n1692), .ip3(n1691), .op(n1694) );
  nor2_1 U818 ( .ip1(n2081), .ip2(n2082), .op(n1792) );
  inv_1 U819 ( .ip(n1498), .op(n796) );
  nor3_1 U820 ( .ip1(n1725), .ip2(n1724), .ip3(n1723), .op(n1726) );
  nor2_1 U821 ( .ip1(n1951), .ip2(n1950), .op(n1952) );
  nor2_1 U822 ( .ip1(n1788), .ip2(n1789), .op(n726) );
  inv_1 U823 ( .ip(n1504), .op(n2065) );
  nand2_1 U824 ( .ip1(n1129), .ip2(n1128), .op(n1208) );
  nor2_1 U825 ( .ip1(n1003), .ip2(n1002), .op(n1004) );
  nand2_1 U826 ( .ip1(n1443), .ip2(n1354), .op(n1446) );
  inv_1 U827 ( .ip(n2028), .op(n712) );
  nor2_1 U828 ( .ip1(n1949), .ip2(n1948), .op(n1950) );
  nand2_1 U829 ( .ip1(n890), .ip2(n889), .op(n1783) );
  nand2_1 U830 ( .ip1(n1637), .ip2(n1636), .op(n2083) );
  nor3_1 U831 ( .ip1(n1955), .ip2(n1943), .ip3(n1947), .op(n1944) );
  nand2_1 U832 ( .ip1(n1612), .ip2(n1611), .op(n2085) );
  nand2_1 U833 ( .ip1(n1025), .ip2(n1024), .op(n1026) );
  and2_1 U834 ( .ip1(n1186), .ip2(n1185), .op(n1722) );
  nand2_1 U835 ( .ip1(n1192), .ip2(n1191), .op(n1678) );
  and2_1 U836 ( .ip1(n1548), .ip2(n1547), .op(n1770) );
  and2_1 U837 ( .ip1(n1554), .ip2(n1553), .op(n1772) );
  nand2_1 U838 ( .ip1(n1089), .ip2(n1088), .op(n1098) );
  nor2_1 U839 ( .ip1(n1188), .ip2(n1187), .op(n1192) );
  xor2_2 U840 ( .ip1(n2046), .ip2(n2045), .op(n1443) );
  nor2_1 U841 ( .ip1(n1550), .ip2(n1549), .op(n1554) );
  nand2_1 U842 ( .ip1(n1125), .ip2(multQ[14]), .op(n1155) );
  nand2_1 U843 ( .ip1(n1599), .ip2(n1598), .op(n2002) );
  nor2_1 U844 ( .ip1(n1606), .ip2(n1605), .op(n1612) );
  nor2_1 U845 ( .ip1(n1610), .ip2(n1609), .op(n1611) );
  nor2_1 U846 ( .ip1(n886), .ip2(n885), .op(n890) );
  nor2_1 U847 ( .ip1(n1629), .ip2(n1628), .op(n1637) );
  nor2_1 U848 ( .ip1(n1635), .ip2(n1634), .op(n1636) );
  nor2_1 U849 ( .ip1(aBQ[0]), .ip2(n2203), .op(n2200) );
  nor2_1 U850 ( .ip1(n1546), .ip2(n1545), .op(n1547) );
  nor2_1 U851 ( .ip1(n888), .ip2(n887), .op(n889) );
  nor2_1 U852 ( .ip1(n1552), .ip2(n1551), .op(n1553) );
  inv_1 U853 ( .ip(n1417), .op(n2006) );
  nor2_1 U854 ( .ip1(n842), .ip2(n841), .op(n848) );
  inv_4 U855 ( .ip(n1342), .op(n714) );
  nand2_1 U856 ( .ip1(n1812), .ip2(n1811), .op(n1088) );
  nor2_1 U857 ( .ip1(n1940), .ip2(n1020), .op(n1030) );
  nor2_1 U858 ( .ip1(n1190), .ip2(n1189), .op(n1191) );
  nor2_1 U859 ( .ip1(aAQ[0]), .ip2(n2219), .op(n2216) );
  mux2_1 U860 ( .ip1(n1965), .ip2(n1964), .s(n1653), .op(n1654) );
  inv_1 U861 ( .ip(n916), .op(n719) );
  inv_1 U862 ( .ip(n1029), .op(n1024) );
  xnor2_1 U863 ( .ip1(n950), .ip2(n949), .op(n951) );
  nor2_1 U864 ( .ip1(n1607), .ip2(n1630), .op(n1610) );
  inv_1 U865 ( .ip(n1660), .op(n1653) );
  nand2_1 U866 ( .ip1(n955), .ip2(n1104), .op(n1047) );
  nor2_2 U867 ( .ip1(n1019), .ip2(n1018), .op(n1945) );
  inv_1 U868 ( .ip(n1340), .op(n1797) );
  nand2_1 U869 ( .ip1(n1819), .ip2(n2096), .op(n2110) );
  nand2_1 U870 ( .ip1(n1090), .ip2(n1091), .op(n1029) );
  buf_1 U871 ( .ip(n1340), .op(n2084) );
  nand2_1 U872 ( .ip1(n1651), .ip2(n1650), .op(n1660) );
  buf_1 U873 ( .ip(n2156), .op(n1273) );
  buf_4 U874 ( .ip(n1285), .op(n716) );
  nor2_1 U875 ( .ip1(n958), .ip2(n1106), .op(n975) );
  inv_1 U876 ( .ip(n1802), .op(n895) );
  inv_1 U877 ( .ip(n1017), .op(n1809) );
  nor2_1 U878 ( .ip1(n2139), .ip2(n2138), .op(n2140) );
  xnor2_1 U879 ( .ip1(counterQ[0]), .ip2(n1437), .op(n1438) );
  nand2_1 U880 ( .ip1(n2224), .ip2(aAQ[3]), .op(n2215) );
  inv_1 U881 ( .ip(n1992), .op(n1406) );
  nor2_2 U882 ( .ip1(n1017), .ip2(n1077), .op(n1018) );
  nand2_1 U883 ( .ip1(n2208), .ip2(aBQ[3]), .op(n2199) );
  nor2_1 U884 ( .ip1(aBQ[4]), .ip2(aBQ[7]), .op(n2197) );
  inv_1 U885 ( .ip(partialQ[13]), .op(n1882) );
  and2_1 U886 ( .ip1(aBQ[1]), .ip2(aBQ[0]), .op(n2208) );
  buf_1 U887 ( .ip(ramBQ[3]), .op(n839) );
  inv_1 U888 ( .ip(ramAQ[2]), .op(n1614) );
  nor2_1 U889 ( .ip1(aBQ[6]), .ip2(aBQ[5]), .op(n2198) );
  inv_1 U890 ( .ip(partialQ[14]), .op(n1154) );
  inv_1 U891 ( .ip(n1463), .op(n717) );
  nor2_1 U892 ( .ip1(aAQ[6]), .ip2(aAQ[5]), .op(n2214) );
  nor2_1 U893 ( .ip1(aAQ[4]), .ip2(aAQ[7]), .op(n2213) );
  and2_1 U894 ( .ip1(aAQ[1]), .ip2(aAQ[0]), .op(n2224) );
  inv_1 U895 ( .ip(partialQ[11]), .op(n1142) );
  inv_1 U896 ( .ip(aBQ[1]), .op(n2204) );
  inv_2 U897 ( .ip(reset), .op(n1303) );
  nor2_2 U898 ( .ip1(n718), .ip2(n756), .op(n757) );
  nand2_1 U899 ( .ip1(n755), .ip2(n754), .op(n718) );
  nand2_1 U900 ( .ip1(n731), .ip2(n730), .op(n729) );
  nand2_1 U901 ( .ip1(n2136), .ip2(n720), .op(n571) );
  nand2_1 U902 ( .ip1(n2123), .ip2(\mult/productQ [22]), .op(n720) );
  nand2_1 U903 ( .ip1(multQ[7]), .ip2(n790), .op(n781) );
  nand2_1 U904 ( .ip1(n765), .ip2(n766), .op(n790) );
  inv_2 U905 ( .ip(n838), .op(n824) );
  nand2_4 U906 ( .ip1(n864), .ip2(n1275), .op(n1727) );
  nand2_1 U907 ( .ip1(n1727), .ip2(\mult/storeQ [11]), .op(n1677) );
  nand3_1 U908 ( .ip1(n724), .ip2(n1802), .ip3(n1793), .op(n723) );
  nand3_2 U909 ( .ip1(n865), .ip2(n896), .ip3(n714), .op(n1529) );
  nor2_1 U910 ( .ip1(counterQ[13]), .ip2(counterQ[9]), .op(n748) );
  nand2_1 U911 ( .ip1(n727), .ip2(n728), .op(n732) );
  nor2_2 U912 ( .ip1(counterQ[3]), .ip2(counterQ[13]), .op(n727) );
  nor2_2 U913 ( .ip1(counterQ[9]), .ip2(counterQ[8]), .op(n728) );
  nor2_2 U914 ( .ip1(n732), .ip2(n729), .op(n765) );
  nor2_2 U915 ( .ip1(counterQ[15]), .ip2(counterQ[4]), .op(n730) );
  nor2_2 U916 ( .ip1(counterQ[14]), .ip2(counterQ[1]), .op(n731) );
  nor2_2 U917 ( .ip1(n761), .ip2(n760), .op(n766) );
  nand2_2 U918 ( .ip1(n733), .ip2(n1456), .op(n760) );
  nor2_2 U919 ( .ip1(counterQ[5]), .ip2(counterQ[7]), .op(n733) );
  inv_2 U920 ( .ip(counterQ[11]), .op(n1456) );
  nand2_2 U921 ( .ip1(n734), .ip2(n735), .op(n761) );
  nor2_2 U922 ( .ip1(counterQ[2]), .ip2(counterQ[10]), .op(n734) );
  nor2_2 U923 ( .ip1(counterQ[6]), .ip2(counterQ[12]), .op(n735) );
  nor2_1 U924 ( .ip1(counterQ[7]), .ip2(counterQ[5]), .op(n759) );
  and2_1 U925 ( .ip1(n1149), .ip2(n1148), .op(n736) );
  inv_2 U926 ( .ip(n736), .op(n1899) );
  nand2_2 U927 ( .ip1(n923), .ip2(n1734), .op(n917) );
  nand2_2 U928 ( .ip1(n861), .ip2(\mult/counterQ [3]), .op(n862) );
  nand3_1 U929 ( .ip1(n1734), .ip2(n1802), .ip3(n714), .op(n899) );
  nor2_1 U930 ( .ip1(n2138), .ip2(n1846), .op(n2129) );
  nand2_1 U931 ( .ip1(n1824), .ip2(n1823), .op(n2141) );
  inv_1 U932 ( .ip(n1151), .op(n2015) );
  inv_1 U933 ( .ip(n1633), .op(n878) );
  inv_1 U934 ( .ip(multQ[2]), .op(n785) );
  inv_1 U935 ( .ip(n1031), .op(n1023) );
  inv_1 U936 ( .ip(n1030), .op(n1025) );
  mux2_1 U937 ( .ip1(n1735), .ip2(n1975), .s(n1734), .op(n2082) );
  inv_2 U938 ( .ip(\mult/counterQ [1]), .op(n1173) );
  inv_1 U939 ( .ip(n1001), .op(n1002) );
  inv_1 U940 ( .ip(n1000), .op(n1003) );
  inv_1 U941 ( .ip(n1649), .op(n1651) );
  inv_1 U942 ( .ip(aBQ[8]), .op(n2195) );
  inv_1 U943 ( .ip(aAQ[8]), .op(n2211) );
  inv_1 U944 ( .ip(n1850), .op(n1845) );
  nand2_1 U945 ( .ip1(n738), .ip2(n1220), .op(n1494) );
  mux2_1 U946 ( .ip1(n1577), .ip2(n1770), .s(\mult/counterQ [2]), .op(n1578)
         );
  inv_1 U947 ( .ip(n1359), .op(n1470) );
  xnor2_1 U948 ( .ip1(n1406), .ip2(n1994), .op(n1995) );
  nor2_1 U949 ( .ip1(n2006), .ip2(n1986), .op(n1987) );
  inv_1 U950 ( .ip(n1249), .op(n1250) );
  inv_1 U951 ( .ip(n2083), .op(n1974) );
  xnor2_1 U952 ( .ip1(n1968), .ip2(n1967), .op(n1969) );
  nor2_1 U953 ( .ip1(n1648), .ip2(n1966), .op(n1967) );
  inv_1 U954 ( .ip(n1772), .op(n1773) );
  nor2_1 U955 ( .ip1(n941), .ip2(n940), .op(n942) );
  nor2_1 U956 ( .ip1(n1680), .ip2(n1679), .op(n1681) );
  inv_1 U957 ( .ip(aAQ[1]), .op(n2220) );
  nand2_1 U958 ( .ip1(n2130), .ip2(n2129), .op(n2131) );
  nor2_1 U959 ( .ip1(n2127), .ip2(n2126), .op(n2132) );
  inv_1 U960 ( .ip(n2107), .op(n2109) );
  xnor2_1 U961 ( .ip1(n979), .ip2(n978), .op(n980) );
  inv_1 U962 ( .ip(n1678), .op(n1565) );
  mux2_1 U963 ( .ip1(n1719), .ip2(n1721), .s(n1734), .op(n1730) );
  mux2_1 U964 ( .ip1(n1686), .ip2(n1540), .s(n1734), .op(n1541) );
  mux2_1 U965 ( .ip1(n1798), .ip2(n2085), .s(\mult/counterQ [2]), .op(n1641)
         );
  nand2_1 U966 ( .ip1(n824), .ip2(n839), .op(n840) );
  nor2_1 U967 ( .ip1(n2017), .ip2(n2015), .op(n1888) );
  nand2_1 U968 ( .ip1(n1125), .ip2(multQ[15]), .op(n1126) );
  nand2_1 U969 ( .ip1(n975), .ip2(n959), .op(n1080) );
  inv_1 U970 ( .ip(n820), .op(n821) );
  nand2_1 U971 ( .ip1(n824), .ip2(ramBQ[7]), .op(n825) );
  nand2_1 U972 ( .ip1(n882), .ip2(n881), .op(n883) );
  nand2_1 U973 ( .ip1(n880), .ip2(n879), .op(n884) );
  inv_1 U974 ( .ip(n1955), .op(n1949) );
  inv_1 U975 ( .ip(n1947), .op(n1948) );
  inv_1 U976 ( .ip(n2129), .op(n1847) );
  nor2_1 U977 ( .ip1(n1184), .ip2(n1183), .op(n1185) );
  nor2_1 U978 ( .ip1(n1175), .ip2(n1174), .op(n1176) );
  nor2_1 U979 ( .ip1(n1544), .ip2(n1543), .op(n1548) );
  inv_1 U980 ( .ip(n1669), .op(n1589) );
  nand2_1 U981 ( .ip1(n1617), .ip2(n1616), .op(n1623) );
  nand2_1 U982 ( .ip1(n1621), .ip2(n1620), .op(n1622) );
  nand2_1 U983 ( .ip1(n1602), .ip2(n1601), .op(n1798) );
  nand2_1 U984 ( .ip1(n2058), .ip2(n2057), .op(n2068) );
  nand3_1 U985 ( .ip1(n1296), .ip2(wrAddr[1]), .ip3(n1298), .op(n1281) );
  nor2_1 U986 ( .ip1(wrAddr[3]), .ip2(wrAddr[2]), .op(n1296) );
  inv_1 U987 ( .ip(wrAddr[0]), .op(n1298) );
  nor2_1 U988 ( .ip1(n2026), .ip2(n2025), .op(n2027) );
  nand2_1 U989 ( .ip1(n712), .ip2(n2024), .op(n2025) );
  nand2_1 U990 ( .ip1(n740), .ip2(n2031), .op(n2033) );
  xnor2_1 U991 ( .ip1(n1413), .ip2(n1411), .op(n1412) );
  xnor2_1 U992 ( .ip1(n1433), .ip2(n1431), .op(n1432) );
  inv_1 U993 ( .ip(n1428), .op(n1429) );
  nand2_1 U994 ( .ip1(n1111), .ip2(n1110), .op(n1112) );
  inv_1 U995 ( .ip(n1881), .op(n1870) );
  nand2_1 U996 ( .ip1(n1060), .ip2(n1059), .op(n1061) );
  nor2_1 U997 ( .ip1(n1033), .ip2(n1032), .op(n1034) );
  nand3_1 U998 ( .ip1(n1028), .ip2(n1027), .ip3(n1026), .op(n1035) );
  nand2_1 U999 ( .ip1(n1023), .ip2(n1024), .op(n1027) );
  nor2_1 U1000 ( .ip1(n1118), .ip2(n961), .op(n949) );
  nor2_1 U1001 ( .ip1(n1005), .ip2(n1004), .op(n1006) );
  mux2_1 U1002 ( .ip1(n1810), .ip2(n1809), .s(n1000), .op(n1005) );
  nand2_1 U1003 ( .ip1(n1655), .ip2(n1654), .op(n1665) );
  nand2_1 U1004 ( .ip1(n1652), .ip2(n1653), .op(n1655) );
  inv_1 U1005 ( .ip(n1661), .op(n1652) );
  nor2_1 U1006 ( .ip1(n1757), .ip2(n1756), .op(n1758) );
  nor3_1 U1007 ( .ip1(wrAddr[1]), .ip2(n1298), .ip3(n1297), .op(n1304) );
  inv_1 U1008 ( .ip(n1995), .op(n1996) );
  xnor2_1 U1009 ( .ip1(n1989), .ip2(n1987), .op(n1988) );
  xnor2_1 U1010 ( .ip1(n1398), .ip2(n2040), .op(n2041) );
  xnor2_1 U1011 ( .ip1(n1401), .ip2(n1418), .op(n1419) );
  nand2_1 U1012 ( .ip1(n1251), .ip2(n1250), .op(n1261) );
  mux2_1 U1013 ( .ip1(n1337), .ip2(n1280), .s(n1802), .op(n630) );
  xnor2_1 U1014 ( .ip1(n1456), .ip2(n1455), .op(n1457) );
  inv_1 U1015 ( .ip(n1969), .op(n1970) );
  xnor2_1 U1016 ( .ip1(n2048), .ip2(n2047), .op(n2050) );
  xnor2_1 U1017 ( .ip1(n943), .ip2(n942), .op(n944) );
  mux2_1 U1018 ( .ip1(n1276), .ip2(n1341), .s(n1734), .op(n628) );
  nand2_1 U1019 ( .ip1(n737), .ip2(n2049), .op(n2001) );
  xnor2_1 U1020 ( .ip1(n1463), .ip2(n1461), .op(n1462) );
  xnor2_1 U1021 ( .ip1(n1449), .ip2(n1447), .op(n1448) );
  xnor2_1 U1022 ( .ip1(n2008), .ip2(n2007), .op(n2009) );
  xnor2_1 U1023 ( .ip1(n1425), .ip2(n1993), .op(n1424) );
  nand2_1 U1024 ( .ip1(n2207), .ip2(aBQ[3]), .op(n2210) );
  and2_1 U1025 ( .ip1(n1292), .ip2(aBQ[4]), .op(n4) );
  and2_1 U1026 ( .ip1(n1292), .ip2(aBQ[5]), .op(n5) );
  and2_1 U1027 ( .ip1(n2161), .ip2(aBQ[6]), .op(n6) );
  and2_1 U1028 ( .ip1(n2161), .ip2(aBQ[7]), .op(n7) );
  nand2_1 U1029 ( .ip1(n2223), .ip2(aAQ[3]), .op(n2227) );
  and2_1 U1030 ( .ip1(n2161), .ip2(aAQ[4]), .op(n12) );
  and2_1 U1031 ( .ip1(n2161), .ip2(aAQ[5]), .op(n13) );
  nand2_1 U1032 ( .ip1(n1857), .ip2(n1856), .op(n1858) );
  xnor2_1 U1033 ( .ip1(n1855), .ip2(n1854), .op(n1857) );
  xnor2_1 U1034 ( .ip1(n2134), .ip2(n2133), .op(n2135) );
  nand2_1 U1035 ( .ip1(n2152), .ip2(n2151), .op(n2153) );
  xnor2_1 U1036 ( .ip1(n2140), .ip2(n2150), .op(n2152) );
  xnor2_1 U1037 ( .ip1(n1828), .ip2(n1827), .op(n1829) );
  nand2_1 U1038 ( .ip1(n2120), .ip2(n2151), .op(n2121) );
  xnor2_1 U1039 ( .ip1(n2119), .ip2(n2118), .op(n2120) );
  xnor2_1 U1040 ( .ip1(n2103), .ip2(n2102), .op(n2104) );
  xnor2_1 U1041 ( .ip1(n1049), .ip2(n1048), .op(n1050) );
  inv_1 U1042 ( .ip(n980), .op(n981) );
  nand2_1 U1043 ( .ip1(n1491), .ip2(n2059), .op(n1493) );
  mux2_1 U1044 ( .ip1(n2049), .ip2(n2064), .s(counterQ[0]), .op(n650) );
  inv_1 U1045 ( .ip(n1216), .op(n1209) );
  and2_1 U1046 ( .ip1(n1178), .ip2(n1973), .op(n738) );
  or2_1 U1047 ( .ip1(n1566), .ip2(n1494), .op(n739) );
  or2_1 U1048 ( .ip1(n2069), .ip2(n712), .op(n740) );
  or2_1 U1049 ( .ip1(n1203), .ip2(n1736), .op(n741) );
  nor2_2 U1050 ( .ip1(n1749), .ip2(n713), .op(n2054) );
  inv_1 U1051 ( .ip(\mult/counterQ [5]), .op(n914) );
  or2_1 U1052 ( .ip1(\mult/storeQ [9]), .ip2(\mult/productQ [9]), .op(n742) );
  or2_1 U1053 ( .ip1(n1908), .ip2(n2069), .op(n743) );
  or2_1 U1054 ( .ip1(n1851), .ip2(n1850), .op(n744) );
  or2_1 U1055 ( .ip1(n2086), .ip2(n1786), .op(n745) );
  or2_1 U1056 ( .ip1(n2115), .ip2(n2114), .op(n746) );
  nor2_2 U1057 ( .ip1(n1282), .ip2(n1311), .op(n1292) );
  inv_1 U1058 ( .ip(n2069), .op(n2024) );
  inv_1 U1059 ( .ip(partialQ[15]), .op(n747) );
  nand2_1 U1061 ( .ip1(n759), .ip2(n1456), .op(n751) );
  nor2_1 U1062 ( .ip1(counterQ[4]), .ip2(counterQ[8]), .op(n749) );
  nand2_1 U1063 ( .ip1(n749), .ip2(n748), .op(n750) );
  nor2_2 U1064 ( .ip1(n750), .ip2(n751), .op(n758) );
  nor2_1 U1065 ( .ip1(counterQ[12]), .ip2(counterQ[10]), .op(n753) );
  nor2_1 U1066 ( .ip1(counterQ[3]), .ip2(counterQ[1]), .op(n755) );
  nor2_1 U1067 ( .ip1(counterQ[14]), .ip2(counterQ[15]), .op(n754) );
  and2_4 U1068 ( .ip1(n757), .ip2(n758), .op(n1146) );
  inv_2 U1069 ( .ip(n1146), .op(n1263) );
  nand2_1 U1070 ( .ip1(n1263), .ip2(multQ[8]), .op(n1163) );
  nand2_1 U1071 ( .ip1(n1163), .ip2(n1700), .op(n1701) );
  nand2_1 U1072 ( .ip1(n766), .ip2(n765), .op(n767) );
  nand2_2 U1073 ( .ip1(multQ[5]), .ip2(n767), .op(n1745) );
  inv_2 U1074 ( .ip(partialQ[5]), .op(n1749) );
  inv_1 U1075 ( .ip(n763), .op(n778) );
  nand2_1 U1076 ( .ip1(multQ[4]), .ip2(n786), .op(n1743) );
  inv_1 U1077 ( .ip(partialQ[4]), .op(n1742) );
  nand2_1 U1078 ( .ip1(n1743), .ip2(n1742), .op(n764) );
  inv_1 U1079 ( .ip(partialQ[7]), .op(n1516) );
  nand2_2 U1080 ( .ip1(n781), .ip2(n1516), .op(n1513) );
  inv_1 U1081 ( .ip(partialQ[6]), .op(n769) );
  nand2_1 U1082 ( .ip1(n767), .ip2(multQ[6]), .op(n768) );
  nand2_2 U1083 ( .ip1(n769), .ip2(n768), .op(n1505) );
  nand2_2 U1084 ( .ip1(n1513), .ip2(n1505), .op(n1236) );
  nor2_2 U1085 ( .ip1(n1236), .ip2(n770), .op(n1863) );
  nand2_1 U1086 ( .ip1(multQ[2]), .ip2(partialQ[2]), .op(n771) );
  nor2_1 U1087 ( .ip1(n1146), .ip2(n771), .op(n1481) );
  inv_1 U1088 ( .ip(n778), .op(n786) );
  nand2_1 U1089 ( .ip1(multQ[3]), .ip2(n786), .op(n773) );
  inv_1 U1090 ( .ip(n773), .op(n774) );
  nand2_2 U1091 ( .ip1(n774), .ip2(partialQ[3]), .op(n1500) );
  nand2_1 U1092 ( .ip1(n1501), .ip2(n1500), .op(n775) );
  nand2_2 U1093 ( .ip1(n1863), .ip2(n775), .op(n1699) );
  nor2_4 U1094 ( .ip1(n1749), .ip2(n1745), .op(n1509) );
  nor2_1 U1095 ( .ip1(multQ[5]), .ip2(partialQ[5]), .op(n776) );
  nand2_1 U1096 ( .ip1(multQ[4]), .ip2(partialQ[4]), .op(n1750) );
  or3_4 U1097 ( .ip1(n1146), .ip2(n776), .ip3(n1750), .op(n1508) );
  inv_4 U1098 ( .ip(n1508), .op(n777) );
  nor2_4 U1099 ( .ip1(n1509), .ip2(n777), .op(n1235) );
  nor2_2 U1100 ( .ip1(n1236), .ip2(n1235), .op(n1862) );
  and2_1 U1101 ( .ip1(partialQ[6]), .ip2(multQ[6]), .op(n779) );
  inv_1 U1102 ( .ip(n778), .op(n1134) );
  nand2_1 U1103 ( .ip1(n779), .ip2(n1134), .op(n780) );
  inv_1 U1104 ( .ip(n780), .op(n1507) );
  nand2_1 U1105 ( .ip1(n1513), .ip2(n1507), .op(n1237) );
  inv_1 U1106 ( .ip(n781), .op(n782) );
  nand2_1 U1107 ( .ip1(n782), .ip2(partialQ[7]), .op(n1514) );
  nand2_2 U1108 ( .ip1(n1237), .ip2(n1514), .op(n1704) );
  nor2_2 U1109 ( .ip1(n1862), .ip2(n1704), .op(n799) );
  inv_1 U1110 ( .ip(multQ[4]), .op(n1225) );
  nand2_1 U1111 ( .ip1(n1225), .ip2(n1742), .op(n783) );
  nand2_1 U1112 ( .ip1(n1227), .ip2(n783), .op(n784) );
  or2_1 U1113 ( .ip1(n784), .ip2(n1236), .op(n798) );
  or2_1 U1114 ( .ip1(n785), .ip2(n1146), .op(n1230) );
  inv_1 U1115 ( .ip(partialQ[2]), .op(n1229) );
  nand2_1 U1116 ( .ip1(n1230), .ip2(n1229), .op(n1487) );
  nand2_1 U1117 ( .ip1(multQ[3]), .ip2(n786), .op(n788) );
  inv_1 U1118 ( .ip(n1231), .op(n789) );
  inv_1 U1119 ( .ip(n789), .op(n1474) );
  nand2_1 U1120 ( .ip1(n1487), .ip2(n1474), .op(n797) );
  nand2_1 U1121 ( .ip1(n790), .ip2(multQ[1]), .op(n794) );
  inv_1 U1122 ( .ip(n794), .op(n791) );
  nand2_2 U1123 ( .ip1(n791), .ip2(partialQ[1]), .op(n1466) );
  nand2_1 U1124 ( .ip1(multQ[0]), .ip2(partialQ[0]), .op(n792) );
  nor2_1 U1125 ( .ip1(n1146), .ip2(n792), .op(n795) );
  inv_1 U1126 ( .ip(partialQ[1]), .op(n793) );
  nand2_1 U1127 ( .ip1(n794), .ip2(n793), .op(n1266) );
  nand2_1 U1128 ( .ip1(n1701), .ip2(n2013), .op(n814) );
  nor2_1 U1129 ( .ip1(n1700), .ip2(n1163), .op(n1243) );
  inv_1 U1130 ( .ip(n1243), .op(n1702) );
  inv_1 U1131 ( .ip(n1702), .op(n806) );
  nor2_1 U1132 ( .ip1(reset), .ip2(state[1]), .op(n800) );
  nand2_2 U1133 ( .ip1(n800), .ip2(state[0]), .op(n805) );
  and2_1 U1134 ( .ip1(partialQ[9]), .ip2(multQ[9]), .op(n801) );
  inv_1 U1135 ( .ip(n1146), .op(n1138) );
  nand2_1 U1136 ( .ip1(n801), .ip2(n1138), .op(n1140) );
  buf_1 U1137 ( .ip(n1140), .op(n1920) );
  nand2_2 U1138 ( .ip1(n1263), .ip2(multQ[9]), .op(n803) );
  inv_1 U1139 ( .ip(partialQ[9]), .op(n802) );
  nand2_4 U1140 ( .ip1(n803), .ip2(n802), .op(n1244) );
  nand2_1 U1141 ( .ip1(n1920), .ip2(n1244), .op(n812) );
  nor3_1 U1142 ( .ip1(n806), .ip2(n2069), .ip3(n812), .op(n804) );
  nand2_1 U1143 ( .ip1(n814), .ip2(n804), .op(n816) );
  nand3_1 U1144 ( .ip1(n812), .ip2(n2024), .ip3(n806), .op(n810) );
  and2_1 U1145 ( .ip1(state[1]), .ip2(n1303), .op(n808) );
  nand2_1 U1146 ( .ip1(n1303), .ip2(n1281), .op(n807) );
  nor2_1 U1147 ( .ip1(n807), .ip2(state[0]), .op(n1301) );
  nor2_2 U1148 ( .ip1(n808), .ip2(n1301), .op(n1917) );
  nand2_1 U1149 ( .ip1(n1293), .ip2(partialQ[9]), .op(n809) );
  nand2_1 U1150 ( .ip1(n812), .ip2(n2059), .op(n813) );
  or2_1 U1151 ( .ip1(n814), .ip2(n813), .op(n815) );
  nand2_4 U1152 ( .ip1(\mult/state [0]), .ip2(n1303), .op(n1295) );
  inv_4 U1153 ( .ip(n1295), .op(n1277) );
  nand2_1 U1154 ( .ip1(\mult/counterQ [5]), .ip2(n1277), .op(n817) );
  and2_1 U1155 ( .ip1(\mult/state [1]), .ip2(n1303), .op(n921) );
  inv_2 U1156 ( .ip(n921), .op(n919) );
  and2_4 U1157 ( .ip1(n817), .ip2(n919), .op(n1275) );
  inv_2 U1158 ( .ip(n1275), .op(n1308) );
  nand2_4 U1159 ( .ip1(n1275), .ip2(n1277), .op(n1342) );
  inv_2 U1160 ( .ip(\mult/counterQ [0]), .op(n1172) );
  buf_1 U1161 ( .ip(n1172), .op(n855) );
  buf_1 U1162 ( .ip(n855), .op(n818) );
  mux2_2 U1163 ( .ip1(n1308), .ip2(n714), .s(n818), .op(n626) );
  buf_1 U1164 ( .ip(\mult/counterQ [1]), .op(n819) );
  nand2_4 U1165 ( .ip1(n1172), .ip2(n819), .op(n866) );
  inv_2 U1166 ( .ip(n866), .op(n1613) );
  inv_2 U1167 ( .ip(n1172), .op(n828) );
  nand2_1 U1168 ( .ip1(n828), .ip2(ramBQ[5]), .op(n820) );
  nand2_1 U1169 ( .ip1(n821), .ip2(n1173), .op(n822) );
  nand2_2 U1170 ( .ip1(n823), .ip2(n822), .op(n932) );
  nand2_1 U1171 ( .ip1(\mult/counterQ [1]), .ip2(\mult/counterQ [0]), .op(n838) );
  nand2_1 U1172 ( .ip1(n1976), .ip2(n825), .op(n826) );
  inv_1 U1173 ( .ip(n826), .op(n931) );
  nand2_2 U1174 ( .ip1(n1618), .ip2(ramBQ[4]), .op(n930) );
  nand2_2 U1175 ( .ip1(n931), .ip2(n930), .op(n893) );
  or2_1 U1176 ( .ip1(n932), .ip2(n893), .op(n865) );
  inv_4 U1177 ( .ip(\mult/counterQ [2]), .op(n1734) );
  inv_1 U1178 ( .ip(ramBQ[12]), .op(n827) );
  or3_1 U1179 ( .ip1(n696), .ip2(n1734), .ip3(n827), .op(n926) );
  and2_1 U1180 ( .ip1(\mult/counterQ [2]), .ip2(ramBQ[13]), .op(n829) );
  nand2_4 U1181 ( .ip1(n1173), .ip2(n828), .op(n869) );
  inv_2 U1182 ( .ip(n869), .op(n1619) );
  nand2_2 U1183 ( .ip1(n829), .ip2(n1619), .op(n925) );
  nand2_1 U1184 ( .ip1(n926), .ip2(n925), .op(n836) );
  nand2_2 U1185 ( .ip1(\mult/counterQ [2]), .ip2(ramBQ[15]), .op(n830) );
  inv_2 U1186 ( .ip(n830), .op(n831) );
  nand2_2 U1187 ( .ip1(n824), .ip2(n831), .op(n832) );
  nand2_2 U1188 ( .ip1(n1976), .ip2(\mult/counterQ [2]), .op(n1340) );
  and2_2 U1189 ( .ip1(n1340), .ip2(n832), .op(n835) );
  and2_1 U1190 ( .ip1(\mult/counterQ [2]), .ip2(ramBQ[14]), .op(n833) );
  nand2_1 U1191 ( .ip1(n833), .ip2(n1613), .op(n834) );
  nand2_2 U1192 ( .ip1(n835), .ip2(n834), .op(n924) );
  or2_2 U1193 ( .ip1(n836), .ip2(n924), .op(n896) );
  nand2_1 U1194 ( .ip1(n865), .ip2(n896), .op(n915) );
  inv_1 U1195 ( .ip(ramBQ[0]), .op(n837) );
  nor2_1 U1196 ( .ip1(n837), .ip2(n696), .op(n842) );
  inv_1 U1197 ( .ip(n838), .op(n877) );
  inv_1 U1198 ( .ip(n840), .op(n841) );
  inv_1 U1199 ( .ip(ramBQ[2]), .op(n843) );
  nor2_1 U1200 ( .ip1(n843), .ip2(n866), .op(n846) );
  inv_1 U1201 ( .ip(ramBQ[1]), .op(n844) );
  nor2_1 U1202 ( .ip1(n844), .ip2(n869), .op(n845) );
  nor2_1 U1203 ( .ip1(n846), .ip2(n845), .op(n847) );
  nand2_1 U1204 ( .ip1(n848), .ip2(n847), .op(n849) );
  nand2_2 U1205 ( .ip1(n849), .ip2(n1976), .op(n863) );
  inv_1 U1206 ( .ip(ramBQ[11]), .op(n850) );
  nand2_1 U1207 ( .ip1(\mult/counterQ [1]), .ip2(\mult/counterQ [0]), .op(
        n1630) );
  nor2_1 U1208 ( .ip1(n850), .ip2(n1630), .op(n853) );
  inv_1 U1209 ( .ip(ramBQ[10]), .op(n851) );
  nor2_1 U1210 ( .ip1(n866), .ip2(n851), .op(n852) );
  nor2_1 U1211 ( .ip1(n853), .ip2(n852), .op(n860) );
  inv_1 U1212 ( .ip(ramBQ[9]), .op(n854) );
  nor2_1 U1213 ( .ip1(n854), .ip2(n869), .op(n858) );
  nand3_1 U1214 ( .ip1(ramBQ[8]), .ip2(n1173), .ip3(n855), .op(n856) );
  inv_1 U1215 ( .ip(n856), .op(n857) );
  nor2_1 U1216 ( .ip1(n858), .ip2(n857), .op(n859) );
  nand2_1 U1217 ( .ip1(n860), .ip2(n859), .op(n861) );
  nand2_4 U1218 ( .ip1(n863), .ip2(n862), .op(n923) );
  nand3_2 U1219 ( .ip1(n915), .ip2(n1277), .ip3(n917), .op(n864) );
  nand2_1 U1220 ( .ip1(n1727), .ip2(\mult/storeQ [23]), .op(n913) );
  inv_1 U1221 ( .ip(n1529), .op(n875) );
  inv_2 U1222 ( .ip(\mult/counterQ [4]), .op(n1802) );
  inv_1 U1223 ( .ip(ramAQ[1]), .op(n1531) );
  buf_1 U1224 ( .ip(n866), .op(n1624) );
  nor2_1 U1225 ( .ip1(n1531), .ip2(n708), .op(n868) );
  inv_1 U1226 ( .ip(ramAQ[3]), .op(n1537) );
  inv_2 U1227 ( .ip(n1618), .op(n1626) );
  nor2_1 U1228 ( .ip1(n1537), .ip2(n1626), .op(n867) );
  inv_1 U1229 ( .ip(ramAQ[0]), .op(n1530) );
  nor2_1 U1230 ( .ip1(n1530), .ip2(n1630), .op(n871) );
  buf_2 U1231 ( .ip(n869), .op(n1632) );
  nor2_1 U1232 ( .ip1(n1614), .ip2(n1632), .op(n870) );
  nor2_1 U1233 ( .ip1(n871), .ip2(n870), .op(n872) );
  nor3_1 U1234 ( .ip1(n1802), .ip2(n2084), .ip3(n2074), .op(n874) );
  nand2_1 U1235 ( .ip1(n875), .ip2(n874), .op(n912) );
  inv_1 U1236 ( .ip(n923), .op(n876) );
  nand2_1 U1237 ( .ip1(n1619), .ip2(ramAQ[10]), .op(n880) );
  inv_1 U1238 ( .ip(ramAQ[8]), .op(n1633) );
  nand2_1 U1239 ( .ip1(n877), .ip2(n878), .op(n879) );
  nand2_1 U1240 ( .ip1(n1618), .ip2(ramAQ[11]), .op(n882) );
  nand2_1 U1241 ( .ip1(n1613), .ip2(ramAQ[9]), .op(n881) );
  nor2_2 U1242 ( .ip1(n884), .ip2(n883), .op(n1669) );
  nand2_1 U1243 ( .ip1(n1669), .ip2(\mult/counterQ [2]), .op(n1790) );
  inv_1 U1244 ( .ip(ramAQ[14]), .op(n1600) );
  nor2_1 U1245 ( .ip1(n1600), .ip2(n1632), .op(n886) );
  inv_1 U1246 ( .ip(ramAQ[15]), .op(n1555) );
  nor2_1 U1247 ( .ip1(n1555), .ip2(n1626), .op(n885) );
  inv_1 U1248 ( .ip(ramAQ[12]), .op(n1608) );
  nor2_1 U1249 ( .ip1(n1608), .ip2(n1630), .op(n888) );
  inv_1 U1250 ( .ip(ramAQ[13]), .op(n1604) );
  nor2_1 U1251 ( .ip1(n1604), .ip2(n708), .op(n887) );
  nand2_1 U1252 ( .ip1(n1783), .ip2(n2081), .op(n891) );
  nand2_1 U1253 ( .ip1(\mult/counterQ [2]), .ip2(\mult/counterQ [3]), .op(
        n1785) );
  nand2_1 U1254 ( .ip1(n891), .ip2(n1785), .op(n892) );
  nand2_1 U1255 ( .ip1(n1790), .ip2(n892), .op(n900) );
  nand3_2 U1256 ( .ip1(n897), .ip2(n714), .ip3(n896), .op(n898) );
  nand2_2 U1257 ( .ip1(n899), .ip2(n898), .op(n1178) );
  inv_2 U1258 ( .ip(n1178), .op(n1219) );
  nor2_1 U1259 ( .ip1(n900), .ip2(n1219), .op(n901) );
  nand2_1 U1260 ( .ip1(n1220), .ip2(n901), .op(n911) );
  nand2_1 U1261 ( .ip1(n1619), .ip2(ramAQ[6]), .op(n903) );
  nand2_1 U1262 ( .ip1(n877), .ip2(ramAQ[4]), .op(n902) );
  nand2_1 U1263 ( .ip1(n903), .ip2(n902), .op(n907) );
  nand2_1 U1264 ( .ip1(n1618), .ip2(ramAQ[7]), .op(n905) );
  nand2_1 U1265 ( .ip1(n1613), .ip2(ramAQ[5]), .op(n904) );
  nand2_1 U1266 ( .ip1(n905), .ip2(n904), .op(n906) );
  nor2_2 U1267 ( .ip1(n907), .ip2(n906), .op(n1786) );
  nand2_1 U1268 ( .ip1(n1734), .ip2(n714), .op(n908) );
  inv_1 U1269 ( .ip(n908), .op(n909) );
  nand2_2 U1270 ( .ip1(n923), .ip2(n909), .op(n1528) );
  inv_1 U1271 ( .ip(n1528), .op(n910) );
  nor2_1 U1272 ( .ip1(\mult/counterQ [2]), .ip2(\mult/counterQ [3]), .op(n1973) );
  and2_1 U1273 ( .ip1(n910), .ip2(n1973), .op(n1170) );
  inv_2 U1274 ( .ip(n1170), .op(n1575) );
  nand4_1 U1275 ( .ip1(n913), .ip2(n912), .ip3(n911), .ip4(n695), .op(n602) );
  nand2_1 U1276 ( .ip1(n1277), .ip2(n914), .op(n916) );
  nand2_2 U1277 ( .ip1(n920), .ip2(n919), .op(n994) );
  inv_1 U1278 ( .ip(n994), .op(n954) );
  inv_1 U1279 ( .ip(n954), .op(n1841) );
  nand2_1 U1280 ( .ip1(n1841), .ip2(\mult/productQ [3]), .op(n946) );
  nor2_1 U1281 ( .ip1(n1295), .ip2(n921), .op(n937) );
  and2_1 U1282 ( .ip1(n1734), .ip2(n937), .op(n922) );
  nand2_2 U1283 ( .ip1(n923), .ip2(n922), .op(n939) );
  inv_1 U1284 ( .ip(n924), .op(n929) );
  nand2_1 U1285 ( .ip1(n926), .ip2(n925), .op(n927) );
  nor2_1 U1286 ( .ip1(n927), .ip2(\mult/counterQ [5]), .op(n928) );
  nand2_1 U1287 ( .ip1(n929), .ip2(n928), .op(n936) );
  and2_1 U1288 ( .ip1(n931), .ip2(n930), .op(n934) );
  nor2_1 U1289 ( .ip1(n932), .ip2(\mult/counterQ [5]), .op(n933) );
  nand2_1 U1290 ( .ip1(n934), .ip2(n933), .op(n935) );
  nand3_2 U1291 ( .ip1(n937), .ip2(n936), .ip3(n935), .op(n938) );
  nand2_4 U1292 ( .ip1(n939), .ip2(n938), .op(n1856) );
  nor2_4 U1293 ( .ip1(\mult/productQ [3]), .ip2(\mult/storeQ [3]), .op(n963)
         );
  and2_1 U1294 ( .ip1(\mult/storeQ [3]), .ip2(\mult/productQ [3]), .op(n966)
         );
  nor2_1 U1295 ( .ip1(n963), .ip2(n966), .op(n943) );
  and2_1 U1296 ( .ip1(\mult/storeQ [2]), .ip2(\mult/productQ [2]), .op(n941)
         );
  nor2_2 U1297 ( .ip1(\mult/storeQ [2]), .ip2(\mult/productQ [2]), .op(n960)
         );
  and2_1 U1298 ( .ip1(\mult/storeQ [1]), .ip2(\mult/productQ [1]), .op(n1118)
         );
  nand2_1 U1299 ( .ip1(\mult/storeQ [0]), .ip2(\mult/productQ [0]), .op(n989)
         );
  nor2_2 U1300 ( .ip1(\mult/storeQ [1]), .ip2(\mult/productQ [1]), .op(n1119)
         );
  nor2_1 U1301 ( .ip1(n989), .ip2(n1119), .op(n961) );
  nor2_1 U1302 ( .ip1(n960), .ip2(n949), .op(n940) );
  nand2_1 U1303 ( .ip1(n1856), .ip2(n944), .op(n945) );
  nand2_1 U1304 ( .ip1(n946), .ip2(n945), .op(n590) );
  buf_1 U1305 ( .ip(\mult/productQ [2]), .op(n947) );
  nand2_1 U1306 ( .ip1(n1841), .ip2(n947), .op(n953) );
  inv_1 U1307 ( .ip(n960), .op(n948) );
  nand2_1 U1308 ( .ip1(\mult/storeQ [2]), .ip2(\mult/productQ [2]), .op(n964)
         );
  and2_1 U1309 ( .ip1(n948), .ip2(n964), .op(n950) );
  nand2_1 U1310 ( .ip1(n1856), .ip2(n951), .op(n952) );
  nand2_1 U1311 ( .ip1(n953), .ip2(n952), .op(n591) );
  inv_1 U1312 ( .ip(n954), .op(n2137) );
  nand2_1 U1313 ( .ip1(n2137), .ip2(\mult/productQ [8]), .op(n973) );
  nor2_2 U1314 ( .ip1(\mult/storeQ [8]), .ip2(\mult/productQ [8]), .op(n1056)
         );
  and2_1 U1315 ( .ip1(\mult/productQ [8]), .ip2(\mult/storeQ [8]), .op(n1058)
         );
  or2_1 U1316 ( .ip1(n1056), .ip2(n1058), .op(n970) );
  or2_1 U1317 ( .ip1(\mult/storeQ [5]), .ip2(\mult/productQ [5]), .op(n1105)
         );
  and2_1 U1318 ( .ip1(\mult/storeQ [4]), .ip2(\mult/productQ [4]), .op(n1109)
         );
  nand2_1 U1319 ( .ip1(n1105), .ip2(n1109), .op(n955) );
  nand2_1 U1320 ( .ip1(\mult/storeQ [5]), .ip2(\mult/productQ [5]), .op(n1104)
         );
  nor2_1 U1321 ( .ip1(\mult/storeQ [7]), .ip2(\mult/productQ [7]), .op(n1041)
         );
  nor2_2 U1322 ( .ip1(\mult/storeQ [6]), .ip2(\mult/productQ [6]), .op(n1043)
         );
  nor2_1 U1323 ( .ip1(n1041), .ip2(n1043), .op(n959) );
  nand2_1 U1324 ( .ip1(n1047), .ip2(n959), .op(n1068) );
  and2_1 U1325 ( .ip1(\mult/storeQ [7]), .ip2(\mult/productQ [7]), .op(n1040)
         );
  nand2_1 U1326 ( .ip1(\mult/productQ [6]), .ip2(\mult/storeQ [6]), .op(n974)
         );
  nor2_1 U1327 ( .ip1(n974), .ip2(n1041), .op(n956) );
  nor2_1 U1328 ( .ip1(n1040), .ip2(n956), .op(n1067) );
  nand2_1 U1329 ( .ip1(n1068), .ip2(n1067), .op(n957) );
  inv_1 U1330 ( .ip(n957), .op(n969) );
  nor2_1 U1331 ( .ip1(\mult/storeQ [5]), .ip2(\mult/productQ [5]), .op(n958)
         );
  nor2_1 U1332 ( .ip1(\mult/storeQ [4]), .ip2(\mult/productQ [4]), .op(n1106)
         );
  inv_1 U1333 ( .ip(n1080), .op(n967) );
  nor2_1 U1334 ( .ip1(n960), .ip2(n963), .op(n962) );
  nand2_1 U1335 ( .ip1(n962), .ip2(n961), .op(n1075) );
  nand2_1 U1336 ( .ip1(n962), .ip2(n1118), .op(n1074) );
  nor2_2 U1337 ( .ip1(n964), .ip2(n963), .op(n965) );
  nor2_2 U1338 ( .ip1(n966), .ip2(n965), .op(n1073) );
  nand3_1 U1339 ( .ip1(n1075), .ip2(n1074), .ip3(n1073), .op(n976) );
  nand2_1 U1340 ( .ip1(n967), .ip2(n976), .op(n968) );
  nand2_2 U1341 ( .ip1(n969), .ip2(n968), .op(n1657) );
  xnor2_2 U1342 ( .ip1(n970), .ip2(n1657), .op(n971) );
  nand2_1 U1343 ( .ip1(n1856), .ip2(n971), .op(n972) );
  nand2_1 U1344 ( .ip1(n973), .ip2(n972), .op(n585) );
  inv_1 U1345 ( .ip(n994), .op(n988) );
  inv_1 U1346 ( .ip(n988), .op(n2123) );
  nand2_1 U1347 ( .ip1(n2123), .ip2(\mult/productQ [6]), .op(n983) );
  inv_1 U1348 ( .ip(n974), .op(n1045) );
  or2_1 U1349 ( .ip1(n1043), .ip2(n1045), .op(n979) );
  nand2_1 U1350 ( .ip1(n976), .ip2(n975), .op(n1042) );
  inv_1 U1351 ( .ip(n1047), .op(n977) );
  and2_1 U1352 ( .ip1(n1042), .ip2(n977), .op(n978) );
  nand2_1 U1353 ( .ip1(n1856), .ip2(n981), .op(n982) );
  nand2_1 U1354 ( .ip1(n983), .ip2(n982), .op(n587) );
  nand2_1 U1355 ( .ip1(n1832), .ip2(\mult/productQ [4]), .op(n987) );
  nor2_1 U1356 ( .ip1(n1106), .ip2(n1109), .op(n984) );
  nand3_1 U1357 ( .ip1(n1075), .ip2(n1074), .ip3(n1073), .op(n1108) );
  xor2_1 U1358 ( .ip1(n984), .ip2(n1108), .op(n985) );
  nand2_1 U1359 ( .ip1(n1856), .ip2(n985), .op(n986) );
  nand2_1 U1360 ( .ip1(n987), .ip2(n986), .op(n589) );
  inv_1 U1361 ( .ip(n988), .op(n1832) );
  nand2_1 U1362 ( .ip1(n1832), .ip2(\mult/productQ [0]), .op(n993) );
  nor2_1 U1363 ( .ip1(\mult/storeQ [0]), .ip2(\mult/productQ [0]), .op(n990)
         );
  inv_1 U1364 ( .ip(n989), .op(n1121) );
  nor2_1 U1365 ( .ip1(n990), .ip2(n1121), .op(n991) );
  nand2_1 U1366 ( .ip1(n1856), .ip2(n991), .op(n992) );
  nand2_1 U1367 ( .ip1(n993), .ip2(n992), .op(n593) );
  inv_1 U1368 ( .ip(n994), .op(n1103) );
  inv_1 U1369 ( .ip(n1103), .op(n1117) );
  nand2_1 U1370 ( .ip1(n1117), .ip2(\mult/productQ [13]), .op(n1012) );
  nor2_4 U1371 ( .ip1(\mult/storeQ [12]), .ip2(\mult/productQ [12]), .op(n1810) );
  nor2_4 U1372 ( .ip1(\mult/storeQ [13]), .ip2(\mult/productQ [13]), .op(n1077) );
  and2_1 U1373 ( .ip1(\mult/productQ [13]), .ip2(\mult/storeQ [13]), .op(n1019) );
  nor2_1 U1374 ( .ip1(n1077), .ip2(n1019), .op(n1000) );
  nor2_2 U1375 ( .ip1(\mult/storeQ [10]), .ip2(\mult/productQ [10]), .op(n1659) );
  nor2_2 U1376 ( .ip1(\mult/storeQ [11]), .ip2(\mult/productQ [11]), .op(n1076) );
  nor2_1 U1377 ( .ip1(n1659), .ip2(n1076), .op(n997) );
  nor2_1 U1378 ( .ip1(\mult/storeQ [9]), .ip2(\mult/productQ [9]), .op(n995)
         );
  nor2_1 U1379 ( .ip1(n995), .ip2(n1056), .op(n1656) );
  nand2_1 U1380 ( .ip1(n997), .ip2(n1656), .op(n1070) );
  inv_1 U1381 ( .ip(n1070), .op(n1021) );
  nand2_2 U1382 ( .ip1(n1657), .ip2(n1021), .op(n1954) );
  nor3_1 U1383 ( .ip1(n1810), .ip2(n1003), .ip3(n1954), .op(n1009) );
  nand2_2 U1384 ( .ip1(\mult/productQ [12]), .ip2(\mult/storeQ [12]), .op(
        n1017) );
  nand2_1 U1385 ( .ip1(n742), .ip2(n1058), .op(n996) );
  nand2_1 U1386 ( .ip1(\mult/productQ [9]), .ip2(\mult/storeQ [9]), .op(n1053)
         );
  nand2_2 U1387 ( .ip1(n996), .ip2(n1053), .op(n1648) );
  nand2_2 U1388 ( .ip1(n1648), .ip2(n997), .op(n1812) );
  and2_1 U1389 ( .ip1(\mult/productQ [11]), .ip2(\mult/storeQ [11]), .op(n1649) );
  nand2_1 U1390 ( .ip1(\mult/productQ [10]), .ip2(\mult/storeQ [10]), .op(
        n1964) );
  nor2_1 U1391 ( .ip1(n1964), .ip2(n1076), .op(n998) );
  nand2_1 U1392 ( .ip1(n1812), .ip2(n1811), .op(n1016) );
  inv_1 U1393 ( .ip(n1810), .op(n1079) );
  and2_1 U1394 ( .ip1(n1016), .ip2(n1079), .op(n1001) );
  nor3_1 U1395 ( .ip1(n1809), .ip2(n1000), .ip3(n1001), .op(n999) );
  nand2_1 U1396 ( .ip1(n999), .ip2(n1954), .op(n1007) );
  nand2_1 U1397 ( .ip1(n1007), .ip2(n1006), .op(n1008) );
  nor2_1 U1398 ( .ip1(n1009), .ip2(n1008), .op(n1010) );
  nand2_1 U1399 ( .ip1(n1010), .ip2(n1856), .op(n1011) );
  nand2_1 U1400 ( .ip1(n1012), .ip2(n1011), .op(n580) );
  nand2_1 U1401 ( .ip1(n1117), .ip2(\mult/productQ [15]), .op(n1039) );
  nor2_1 U1402 ( .ip1(\mult/storeQ [15]), .ip2(\mult/productQ [15]), .op(n1069) );
  inv_1 U1403 ( .ip(n1069), .op(n1090) );
  nand2_1 U1404 ( .ip1(\mult/productQ [15]), .ip2(\mult/storeQ [15]), .op(
        n1091) );
  nor2_2 U1405 ( .ip1(n1810), .ip2(n1077), .op(n1956) );
  nor2_2 U1406 ( .ip1(\mult/storeQ [14]), .ip2(\mult/productQ [14]), .op(n1941) );
  inv_1 U1407 ( .ip(n1941), .op(n1013) );
  and2_1 U1408 ( .ip1(n1956), .ip2(n1013), .op(n1015) );
  and2_1 U1409 ( .ip1(n1657), .ip2(n1015), .op(n1032) );
  inv_1 U1410 ( .ip(n1032), .op(n1014) );
  nor3_1 U1411 ( .ip1(n1070), .ip2(n1029), .ip3(n1014), .op(n1036) );
  nand2_1 U1412 ( .ip1(n1016), .ip2(n1015), .op(n1031) );
  and2_1 U1413 ( .ip1(\mult/productQ [14]), .ip2(\mult/storeQ [14]), .op(n1940) );
  nor2_1 U1414 ( .ip1(n1941), .ip2(n1945), .op(n1020) );
  nor2_1 U1415 ( .ip1(n1024), .ip2(n1021), .op(n1022) );
  nand3_1 U1416 ( .ip1(n1031), .ip2(n1030), .ip3(n1022), .op(n1028) );
  nand3_1 U1417 ( .ip1(n1031), .ip2(n1030), .ip3(n1029), .op(n1033) );
  nor3_1 U1418 ( .ip1(n1036), .ip2(n1035), .ip3(n1034), .op(n1037) );
  nand2_1 U1419 ( .ip1(n1037), .ip2(n1856), .op(n1038) );
  nand2_1 U1420 ( .ip1(n1039), .ip2(n1038), .op(n578) );
  nand2_1 U1421 ( .ip1(n1117), .ip2(\mult/productQ [7]), .op(n1052) );
  nor2_1 U1422 ( .ip1(n1041), .ip2(n1040), .op(n1049) );
  inv_1 U1423 ( .ip(n1043), .op(n1046) );
  nor2_1 U1424 ( .ip1(n1043), .ip2(n1042), .op(n1044) );
  not_ab_or_c_or_d U1425 ( .ip1(n1047), .ip2(n1046), .ip3(n1045), .ip4(n1044), 
        .op(n1048) );
  nand2_1 U1426 ( .ip1(n1050), .ip2(n1856), .op(n1051) );
  nand2_1 U1427 ( .ip1(n1052), .ip2(n1051), .op(n586) );
  nand2_1 U1428 ( .ip1(n1841), .ip2(\mult/productQ [9]), .op(n1065) );
  nor2_1 U1429 ( .ip1(\mult/storeQ [9]), .ip2(\mult/productQ [9]), .op(n1055)
         );
  inv_1 U1430 ( .ip(n1053), .op(n1054) );
  nor2_1 U1431 ( .ip1(n1055), .ip2(n1054), .op(n1062) );
  inv_1 U1432 ( .ip(n1056), .op(n1057) );
  nand2_1 U1433 ( .ip1(n1657), .ip2(n1057), .op(n1060) );
  inv_1 U1434 ( .ip(n1058), .op(n1059) );
  xor2_1 U1435 ( .ip1(n1062), .ip2(n1061), .op(n1063) );
  nand2_4 U1436 ( .ip1(n1063), .ip2(n2151), .op(n1064) );
  nand2_1 U1437 ( .ip1(n1065), .ip2(n1064), .op(n584) );
  nand2_1 U1438 ( .ip1(n1808), .ip2(\mult/productQ [16]), .op(n1102) );
  and2_1 U1439 ( .ip1(\mult/productQ [16]), .ip2(\mult/storeQ [16]), .op(n2101) );
  inv_1 U1440 ( .ip(n2101), .op(n1066) );
  or2_1 U1441 ( .ip1(\mult/storeQ [16]), .ip2(\mult/productQ [16]), .op(n2098)
         );
  nand2_1 U1442 ( .ip1(n1066), .ip2(n2098), .op(n1099) );
  nand2_1 U1443 ( .ip1(n1068), .ip2(n1067), .op(n1072) );
  nor2_2 U1444 ( .ip1(n1941), .ip2(n1069), .op(n1093) );
  nand2_1 U1445 ( .ip1(n1093), .ip2(n1956), .op(n1087) );
  nor2_1 U1446 ( .ip1(n1087), .ip2(n1070), .op(n1071) );
  nand2_1 U1447 ( .ip1(n1072), .ip2(n1071), .op(n1086) );
  nand3_1 U1448 ( .ip1(n1075), .ip2(n1074), .ip3(n1073), .op(n1084) );
  nand2_1 U1449 ( .ip1(n1093), .ip2(n1656), .op(n1082) );
  inv_1 U1450 ( .ip(n1659), .op(n1965) );
  inv_1 U1451 ( .ip(n1076), .op(n1650) );
  inv_1 U1452 ( .ip(n1077), .op(n1078) );
  nand4_1 U1453 ( .ip1(n1965), .ip2(n1650), .ip3(n1079), .ip4(n1078), .op(
        n1081) );
  nand2_1 U1454 ( .ip1(n1084), .ip2(n1083), .op(n1085) );
  nand2_2 U1455 ( .ip1(n1086), .ip2(n1085), .op(n1834) );
  inv_1 U1456 ( .ip(n1087), .op(n1089) );
  nand2_1 U1457 ( .ip1(n1090), .ip2(n1940), .op(n1092) );
  nand2_1 U1458 ( .ip1(n1092), .ip2(n1091), .op(n1096) );
  inv_1 U1459 ( .ip(n1093), .op(n1094) );
  nor2_2 U1460 ( .ip1(n1094), .ip2(n1945), .op(n1095) );
  nor2_2 U1461 ( .ip1(n1096), .ip2(n1095), .op(n1097) );
  nand2_2 U1462 ( .ip1(n1098), .ip2(n1097), .op(n1833) );
  nor2_2 U1463 ( .ip1(n1834), .ip2(n1833), .op(n2126) );
  xnor2_2 U1464 ( .ip1(n1099), .ip2(n2126), .op(n1100) );
  inv_1 U1465 ( .ip(n1856), .op(n1960) );
  or2_1 U1466 ( .ip1(n1100), .ip2(n1960), .op(n1101) );
  nand2_1 U1467 ( .ip1(n1102), .ip2(n1101), .op(n577) );
  inv_1 U1468 ( .ip(n1103), .op(n1808) );
  nand2_1 U1469 ( .ip1(n1808), .ip2(\mult/productQ [5]), .op(n1116) );
  and2_1 U1470 ( .ip1(n1105), .ip2(n1104), .op(n1113) );
  inv_1 U1471 ( .ip(n1106), .op(n1107) );
  nand2_1 U1472 ( .ip1(n1108), .ip2(n1107), .op(n1111) );
  inv_1 U1473 ( .ip(n1109), .op(n1110) );
  xor2_1 U1474 ( .ip1(n1113), .ip2(n1112), .op(n1114) );
  nand2_4 U1475 ( .ip1(n2151), .ip2(n1114), .op(n1115) );
  nand2_1 U1476 ( .ip1(n1116), .ip2(n1115), .op(n588) );
  nand2_1 U1477 ( .ip1(n1117), .ip2(\mult/productQ [1]), .op(n1124) );
  nor2_1 U1478 ( .ip1(n1119), .ip2(n1118), .op(n1120) );
  xor2_1 U1479 ( .ip1(n1121), .ip2(n1120), .op(n1122) );
  nand2_4 U1480 ( .ip1(n2151), .ip2(n1122), .op(n1123) );
  nand2_1 U1481 ( .ip1(n1124), .ip2(n1123), .op(n592) );
  inv_1 U1482 ( .ip(n1146), .op(n1125) );
  nand2_1 U1483 ( .ip1(n1126), .ip2(n747), .op(n1129) );
  inv_1 U1484 ( .ip(n1126), .op(n1127) );
  nand2_1 U1485 ( .ip1(n1127), .ip2(partialQ[15]), .op(n1128) );
  inv_1 U1486 ( .ip(n1208), .op(n1130) );
  nand2_1 U1487 ( .ip1(n1130), .ip2(n1354), .op(n1162) );
  and2_1 U1488 ( .ip1(partialQ[10]), .ip2(multQ[10]), .op(n1131) );
  nand2_1 U1489 ( .ip1(n1131), .ip2(n1138), .op(n1132) );
  nand2_1 U1490 ( .ip1(multQ[11]), .ip2(n1134), .op(n1133) );
  nand2_2 U1491 ( .ip1(n1133), .ip2(n1142), .op(n1871) );
  nand2_1 U1492 ( .ip1(n1871), .ip2(n1872), .op(n1136) );
  nand2_1 U1493 ( .ip1(multQ[11]), .ip2(n1134), .op(n1143) );
  inv_1 U1494 ( .ip(n1143), .op(n1135) );
  nand2_1 U1495 ( .ip1(n1136), .ip2(n1873), .op(n1137) );
  inv_1 U1496 ( .ip(n1137), .op(n1898) );
  nand3_1 U1497 ( .ip1(multQ[8]), .ip2(n1138), .ip3(partialQ[8]), .op(n1139)
         );
  nand2_1 U1498 ( .ip1(n1139), .ip2(n1140), .op(n1141) );
  nand2_1 U1499 ( .ip1(n1141), .ip2(n1244), .op(n1877) );
  nand2_1 U1500 ( .ip1(n1143), .ip2(n1142), .op(n1145) );
  nand2_1 U1501 ( .ip1(n1134), .ip2(multQ[10]), .op(n1239) );
  or2_1 U1502 ( .ip1(n1877), .ip2(n1876), .op(n1897) );
  nand2_1 U1503 ( .ip1(n1898), .ip2(n1897), .op(n1207) );
  inv_1 U1504 ( .ip(n1146), .op(n1147) );
  nand2_1 U1505 ( .ip1(multQ[13]), .ip2(n1147), .op(n1156) );
  nand2_1 U1506 ( .ip1(n1156), .ip2(n1882), .op(n1151) );
  nand2_1 U1507 ( .ip1(n1147), .ip2(multQ[12]), .op(n1149) );
  inv_1 U1508 ( .ip(partialQ[12]), .op(n1148) );
  nor2_2 U1509 ( .ip1(n2015), .ip2(n736), .op(n2020) );
  nand2_2 U1510 ( .ip1(n1155), .ip2(n1154), .op(n2023) );
  nand2_2 U1511 ( .ip1(n2020), .ip2(n2023), .op(n1166) );
  inv_2 U1512 ( .ip(n1166), .op(n1206) );
  nand2_1 U1513 ( .ip1(n1207), .ip2(n1206), .op(n1160) );
  inv_1 U1514 ( .ip(n1149), .op(n1150) );
  inv_1 U1515 ( .ip(n1151), .op(n1152) );
  nand2_1 U1516 ( .ip1(n1153), .ip2(n2023), .op(n1158) );
  or2_1 U1517 ( .ip1(n1155), .ip2(n1154), .op(n2022) );
  nor2_1 U1518 ( .ip1(n1882), .ip2(n1156), .op(n2017) );
  nand2_1 U1519 ( .ip1(n2023), .ip2(n2017), .op(n1157) );
  nor2_1 U1520 ( .ip1(n1162), .ip2(n1161), .op(n1168) );
  buf_1 U1521 ( .ip(n1876), .op(n1165) );
  nand2_1 U1522 ( .ip1(n1163), .ip2(n1700), .op(n1164) );
  nand2_1 U1523 ( .ip1(n1164), .ip2(n1244), .op(n1929) );
  nor2_2 U1524 ( .ip1(n1165), .ip2(n1929), .op(n2012) );
  inv_1 U1525 ( .ip(n2012), .op(n1905) );
  nor2_1 U1526 ( .ip1(n1166), .ip2(n1905), .op(n1167) );
  nand2_1 U1527 ( .ip1(n2013), .ip2(n1167), .op(n1215) );
  nand2_1 U1528 ( .ip1(n1168), .ip2(n1215), .op(n1169) );
  inv_1 U1529 ( .ip(n1169), .op(n2159) );
  nand2_1 U1530 ( .ip1(n1618), .ip2(ramAQ[0]), .op(n1719) );
  nor2_1 U1531 ( .ip1(n1802), .ip2(n1719), .op(n1171) );
  nand2_1 U1532 ( .ip1(n1171), .ip2(n1170), .op(n1179) );
  nand2_1 U1533 ( .ip1(n1604), .ip2(n877), .op(n1177) );
  nor2_1 U1534 ( .ip1(n828), .ip2(ramAQ[14]), .op(n1175) );
  nor2_1 U1535 ( .ip1(ramAQ[15]), .ip2(n819), .op(n1174) );
  nand3_1 U1536 ( .ip1(n1177), .ip2(n1176), .ip3(n1626), .op(n1566) );
  nand2_1 U1537 ( .ip1(n1179), .ip2(n739), .op(n1180) );
  inv_1 U1538 ( .ip(n1180), .op(n1205) );
  nor2_1 U1539 ( .ip1(\mult/counterQ [2]), .ip2(n1976), .op(n1796) );
  nor2_1 U1540 ( .ip1(ramAQ[7]), .ip2(n1632), .op(n1182) );
  nor2_1 U1541 ( .ip1(ramAQ[8]), .ip2(n1626), .op(n1181) );
  nor2_1 U1542 ( .ip1(n1182), .ip2(n1181), .op(n1186) );
  nor2_1 U1543 ( .ip1(ramAQ[5]), .ip2(n1630), .op(n1184) );
  nor2_1 U1544 ( .ip1(ramAQ[6]), .ip2(n708), .op(n1183) );
  nor2_1 U1545 ( .ip1(ramAQ[11]), .ip2(n1632), .op(n1188) );
  nor2_1 U1546 ( .ip1(ramAQ[12]), .ip2(n1626), .op(n1187) );
  inv_1 U1547 ( .ip(ramAQ[9]), .op(n1627) );
  and2_1 U1548 ( .ip1(n877), .ip2(n1627), .op(n1190) );
  nor2_1 U1549 ( .ip1(ramAQ[10]), .ip2(n708), .op(n1189) );
  nor2_1 U1550 ( .ip1(n2084), .ip2(n1678), .op(n1200) );
  nor2_1 U1551 ( .ip1(ramAQ[3]), .ip2(n1632), .op(n1194) );
  nor2_1 U1552 ( .ip1(ramAQ[4]), .ip2(n1626), .op(n1193) );
  nor2_1 U1553 ( .ip1(n1194), .ip2(n1193), .op(n1198) );
  and2_1 U1554 ( .ip1(n877), .ip2(n1531), .op(n1196) );
  nor2_1 U1555 ( .ip1(ramAQ[2]), .ip2(n1624), .op(n1195) );
  nor2_1 U1556 ( .ip1(n1196), .ip2(n1195), .op(n1197) );
  nand2_1 U1557 ( .ip1(n1197), .ip2(n1198), .op(n1721) );
  nor2_1 U1558 ( .ip1(n1785), .ip2(n1721), .op(n1199) );
  not_ab_or_c_or_d U1559 ( .ip1(n1796), .ip2(n1722), .ip3(n1200), .ip4(n1199), 
        .op(n1202) );
  or2_1 U1560 ( .ip1(n1202), .ip2(n1795), .op(n1204) );
  inv_1 U1561 ( .ip(\mult/storeQ [16]), .op(n1203) );
  nand3_1 U1562 ( .ip1(n1205), .ip2(n1204), .ip3(n741), .op(n609) );
  nand2_1 U1563 ( .ip1(n1207), .ip2(n1206), .op(n1210) );
  or2_1 U1564 ( .ip1(n1210), .ip2(n1216), .op(n1214) );
  nand2_1 U1565 ( .ip1(n1209), .ip2(n1211), .op(n1213) );
  nand2_1 U1566 ( .ip1(n1293), .ip2(partialQ[15]), .op(n1212) );
  nand3_1 U1567 ( .ip1(n1214), .ip2(n1213), .ip3(n1212), .op(n1218) );
  nor2_1 U1568 ( .ip1(n1216), .ip2(n1215), .op(n1217) );
  nor2_1 U1569 ( .ip1(n1218), .ip2(n1217), .op(n2160) );
  nand2_1 U1570 ( .ip1(n1727), .ip2(\mult/storeQ [7]), .op(n1224) );
  nand2_1 U1571 ( .ip1(n1201), .ip2(n1220), .op(n1576) );
  inv_1 U1572 ( .ip(n1576), .op(n1675) );
  nor2_1 U1573 ( .ip1(n2084), .ip2(n2074), .op(n1221) );
  nand2_1 U1574 ( .ip1(n1675), .ip2(n1221), .op(n1223) );
  inv_1 U1575 ( .ip(n1973), .op(n2086) );
  or2_1 U1576 ( .ip1(n1795), .ip2(n745), .op(n1222) );
  nand3_1 U1577 ( .ip1(n1224), .ip2(n1223), .ip3(n1222), .op(n618) );
  nand2_1 U1578 ( .ip1(n1225), .ip2(n1742), .op(n1226) );
  or2_1 U1579 ( .ip1(n1504), .ip2(n1236), .op(n1866) );
  nand2_1 U1580 ( .ip1(n1466), .ip2(n1228), .op(n1234) );
  nand2_1 U1581 ( .ip1(n1230), .ip2(n1229), .op(n1232) );
  or2_1 U1582 ( .ip1(n1866), .ip2(n1865), .op(n1904) );
  nor2_2 U1583 ( .ip1(n1235), .ip2(n1236), .op(n1703) );
  nand2_1 U1584 ( .ip1(n1237), .ip2(n1514), .op(n1861) );
  nor2_1 U1585 ( .ip1(n1703), .ip2(n1861), .op(n1238) );
  nand3_1 U1586 ( .ip1(n1904), .ip2(n1699), .ip3(n1238), .op(n1242) );
  nor2_1 U1587 ( .ip1(n1922), .ip2(n1929), .op(n1241) );
  nand2_1 U1588 ( .ip1(n1871), .ip2(n1873), .op(n1247) );
  nand2_1 U1589 ( .ip1(n1247), .ip2(n1354), .op(n1254) );
  and2_1 U1590 ( .ip1(n1241), .ip2(n1255), .op(n1240) );
  nand2_1 U1591 ( .ip1(n1242), .ip2(n1240), .op(n1262) );
  nand2_1 U1592 ( .ip1(n1242), .ip2(n1241), .op(n1251) );
  inv_1 U1593 ( .ip(n1922), .op(n1246) );
  nand2_1 U1594 ( .ip1(n1243), .ip2(n1244), .op(n1919) );
  nand2_1 U1595 ( .ip1(n1920), .ip2(n1919), .op(n1245) );
  nand2_1 U1596 ( .ip1(n1246), .ip2(n1245), .op(n1253) );
  inv_1 U1597 ( .ip(n1872), .op(n1252) );
  inv_1 U1598 ( .ip(n1252), .op(n1921) );
  nor3_1 U1599 ( .ip1(n1921), .ip2(n2069), .ip3(n1247), .op(n1248) );
  nand2_1 U1600 ( .ip1(n1253), .ip2(n1248), .op(n1249) );
  nand2_1 U1601 ( .ip1(n1253), .ip2(n1252), .op(n1256) );
  inv_1 U1602 ( .ip(n1254), .op(n1255) );
  nand2_1 U1603 ( .ip1(n1256), .ip2(n1255), .op(n1258) );
  nand2_1 U1604 ( .ip1(n1293), .ip2(partialQ[11]), .op(n1257) );
  nand2_1 U1605 ( .ip1(n1258), .ip2(n1257), .op(n1259) );
  inv_1 U1606 ( .ip(n1259), .op(n1260) );
  nand3_1 U1607 ( .ip1(n1262), .ip2(n1261), .ip3(n1260), .op(n534) );
  inv_1 U1608 ( .ip(multQ[0]), .op(n1265) );
  inv_1 U1609 ( .ip(n1263), .op(n1264) );
  nor2_2 U1610 ( .ip1(n1265), .ip2(n1264), .op(n1359) );
  inv_1 U1611 ( .ip(partialQ[0]), .op(n1467) );
  or2_1 U1612 ( .ip1(n1470), .ip2(n1467), .op(n1361) );
  inv_1 U1613 ( .ip(n1266), .op(n1468) );
  inv_1 U1614 ( .ip(n1468), .op(n1267) );
  nand2_1 U1615 ( .ip1(n1466), .ip2(n1267), .op(n1268) );
  xor2_1 U1616 ( .ip1(n1361), .ip2(n1268), .op(n1269) );
  nand2_4 U1617 ( .ip1(n1269), .ip2(n2059), .op(n1271) );
  nand2_1 U1618 ( .ip1(n1293), .ip2(partialQ[1]), .op(n1270) );
  inv_1 U1619 ( .ip(\mult/state [1]), .op(n1272) );
  nor2_1 U1620 ( .ip1(\mult/state [0]), .ip2(n1272), .op(n2156) );
  nand2_2 U1621 ( .ip1(state[0]), .ip2(state[1]), .op(n529) );
  nor2_2 U1622 ( .ip1(reset), .ip2(n529), .op(n1285) );
  nand2_1 U1623 ( .ip1(n1630), .ip2(n1277), .op(n1274) );
  and2_1 U1624 ( .ip1(n1275), .ip2(n1274), .op(n1343) );
  inv_1 U1625 ( .ip(n1343), .op(n1276) );
  nand2_1 U1626 ( .ip1(n877), .ip2(n714), .op(n1279) );
  inv_1 U1627 ( .ip(n1279), .op(n1341) );
  nand2_1 U1628 ( .ip1(n1277), .ip2(n1785), .op(n1278) );
  nand2_1 U1629 ( .ip1(n1343), .ip2(n1278), .op(n1337) );
  nor2_1 U1630 ( .ip1(n1785), .ip2(n1279), .op(n1280) );
  nand2_1 U1631 ( .ip1(n2210), .ip2(n2209), .op(n3) );
  nand2_1 U1632 ( .ip1(n2227), .ip2(n2226), .op(n11) );
  nor3_1 U1633 ( .ip1(n1281), .ip2(state[1]), .ip3(state[0]), .op(n1282) );
  nand2_2 U1634 ( .ip1(n529), .ip2(n1303), .op(n1311) );
  buf_2 U1635 ( .ip(n1292), .op(n2161) );
  nand2_1 U1636 ( .ip1(n2212), .ip2(n2211), .op(n1284) );
  nand2_1 U1637 ( .ip1(n2214), .ip2(n2213), .op(n1283) );
  nor2_1 U1638 ( .ip1(n1284), .ip2(n1283), .op(n1286) );
  nand3_2 U1639 ( .ip1(n1286), .ip2(n716), .ip3(n2215), .op(n2219) );
  inv_1 U1640 ( .ip(n2219), .op(n2225) );
  nand2_1 U1641 ( .ip1(n2225), .ip2(n2220), .op(n1287) );
  nand2_1 U1642 ( .ip1(n2221), .ip2(n1287), .op(n2223) );
  nand2_1 U1643 ( .ip1(n2196), .ip2(n2195), .op(n1289) );
  nand2_1 U1644 ( .ip1(n2198), .ip2(n2197), .op(n1288) );
  nor2_1 U1645 ( .ip1(n1289), .ip2(n1288), .op(n1290) );
  nand3_2 U1646 ( .ip1(n1290), .ip2(n716), .ip3(n2199), .op(n2203) );
  inv_1 U1647 ( .ip(n2203), .op(n2228) );
  nand2_1 U1648 ( .ip1(n2228), .ip2(n2204), .op(n1291) );
  nand2_1 U1649 ( .ip1(n2205), .ip2(n1291), .op(n2207) );
  inv_1 U1650 ( .ip(n2202), .op(n1) );
  inv_1 U1651 ( .ip(n2218), .op(n9) );
  buf_4 U1652 ( .ip(n1293), .op(n2064) );
  inv_1 U1653 ( .ip(state[1]), .op(n1305) );
  nor2_1 U1654 ( .ip1(state[0]), .ip2(n1305), .op(n2232) );
  nor2_1 U1655 ( .ip1(\mult/state [1]), .ip2(\mult/counterQ [5]), .op(n1294)
         );
  nor2_1 U1656 ( .ip1(n1295), .ip2(n1294), .op(n634) );
  inv_1 U1657 ( .ip(state[0]), .op(n1299) );
  inv_1 U1658 ( .ip(n1296), .op(n1297) );
  nand3_1 U1659 ( .ip1(n1299), .ip2(n1304), .ip3(n1305), .op(n528) );
  nor2_1 U1660 ( .ip1(n1304), .ip2(state[1]), .op(n1300) );
  nand2_1 U1661 ( .ip1(n1301), .ip2(n1300), .op(n1302) );
  and2_1 U1662 ( .ip1(n1302), .ip2(n1303), .op(n2162) );
  nand3_1 U1663 ( .ip1(n1305), .ip2(n1304), .ip3(n1303), .op(n1306) );
  nand2_1 U1664 ( .ip1(n2069), .ip2(n1306), .op(n683) );
  nand2_1 U1665 ( .ip1(n1632), .ip2(n708), .op(n1307) );
  nand2_1 U1666 ( .ip1(n714), .ip2(n1307), .op(n1310) );
  nand2_1 U1667 ( .ip1(n1308), .ip2(n819), .op(n1309) );
  nand2_1 U1668 ( .ip1(n1310), .ip2(n1309), .op(n627) );
  nand2_1 U1669 ( .ip1(n1387), .ip2(ramAQ[8]), .op(n1312) );
  nand2_1 U1670 ( .ip1(n1312), .ip2(n2186), .op(n675) );
  nand2_1 U1671 ( .ip1(n1387), .ip2(ramAQ[6]), .op(n1313) );
  nand2_1 U1672 ( .ip1(n1313), .ip2(n2185), .op(n673) );
  nand2_1 U1673 ( .ip1(n1387), .ip2(ramAQ[5]), .op(n1314) );
  nand2_1 U1674 ( .ip1(n1314), .ip2(n2184), .op(n672) );
  nand2_1 U1675 ( .ip1(n1387), .ip2(ramBQ[7]), .op(n1315) );
  nand2_1 U1676 ( .ip1(n1315), .ip2(n2170), .op(n658) );
  nand2_1 U1677 ( .ip1(n1387), .ip2(ramAQ[2]), .op(n1316) );
  nand2_1 U1678 ( .ip1(n1316), .ip2(n2180), .op(n669) );
  nand2_1 U1679 ( .ip1(n1387), .ip2(ramAQ[1]), .op(n1317) );
  nand2_1 U1680 ( .ip1(n1317), .ip2(n2181), .op(n668) );
  nand2_1 U1681 ( .ip1(n1387), .ip2(ramAQ[3]), .op(n1318) );
  nand2_1 U1682 ( .ip1(n1318), .ip2(n2183), .op(n670) );
  nand2_1 U1683 ( .ip1(n1387), .ip2(ramAQ[4]), .op(n1319) );
  nand2_1 U1684 ( .ip1(n1319), .ip2(n2182), .op(n671) );
  nand2_1 U1685 ( .ip1(n1387), .ip2(ramBQ[8]), .op(n1320) );
  nand2_1 U1686 ( .ip1(n1320), .ip2(n2177), .op(n659) );
  nand2_1 U1687 ( .ip1(n1387), .ip2(ramBQ[15]), .op(n1321) );
  nand2_1 U1688 ( .ip1(n1321), .ip2(n2164), .op(n666) );
  nand2_1 U1689 ( .ip1(n1387), .ip2(ramBQ[14]), .op(n1322) );
  nand2_1 U1690 ( .ip1(n1322), .ip2(n2166), .op(n665) );
  nand2_1 U1691 ( .ip1(n1387), .ip2(ramBQ[3]), .op(n1323) );
  nand2_1 U1692 ( .ip1(n1323), .ip2(n2171), .op(n654) );
  nand2_1 U1693 ( .ip1(n1387), .ip2(ramBQ[2]), .op(n1324) );
  nand2_1 U1694 ( .ip1(n1324), .ip2(n2173), .op(n653) );
  nand2_1 U1695 ( .ip1(n1387), .ip2(ramBQ[1]), .op(n1325) );
  nand2_1 U1696 ( .ip1(n1325), .ip2(n2174), .op(n652) );
  nand2_1 U1697 ( .ip1(n1387), .ip2(ramBQ[11]), .op(n1326) );
  nand2_1 U1698 ( .ip1(n1326), .ip2(n2175), .op(n662) );
  nand2_1 U1699 ( .ip1(n1387), .ip2(ramBQ[13]), .op(n1327) );
  nand2_1 U1700 ( .ip1(n1327), .ip2(n2165), .op(n664) );
  nand2_1 U1701 ( .ip1(n1387), .ip2(ramBQ[9]), .op(n1328) );
  nand2_1 U1702 ( .ip1(n1328), .ip2(n2178), .op(n660) );
  nand2_1 U1703 ( .ip1(n1387), .ip2(ramBQ[10]), .op(n1329) );
  nand2_1 U1704 ( .ip1(n1329), .ip2(n2176), .op(n661) );
  nand2_1 U1705 ( .ip1(n1387), .ip2(ramBQ[0]), .op(n1330) );
  nand2_1 U1706 ( .ip1(n1330), .ip2(n2172), .op(n651) );
  nand2_1 U1707 ( .ip1(n1387), .ip2(ramBQ[5]), .op(n1331) );
  nand2_1 U1708 ( .ip1(n1331), .ip2(n2169), .op(n656) );
  nand2_1 U1709 ( .ip1(n1387), .ip2(ramBQ[4]), .op(n1332) );
  nand2_1 U1710 ( .ip1(n1332), .ip2(n2167), .op(n655) );
  nand2_1 U1711 ( .ip1(n1387), .ip2(ramBQ[6]), .op(n1333) );
  nand2_1 U1712 ( .ip1(n1333), .ip2(n2168), .op(n657) );
  nand2_1 U1713 ( .ip1(n1387), .ip2(ramBQ[12]), .op(n1334) );
  nand2_1 U1714 ( .ip1(n1334), .ip2(n2163), .op(n663) );
  nand2_1 U1715 ( .ip1(n1387), .ip2(ramAQ[0]), .op(n1335) );
  nand2_1 U1716 ( .ip1(n1335), .ip2(n2179), .op(n667) );
  nor2_1 U1717 ( .ip1(n1802), .ip2(n1785), .op(n1336) );
  nand2_1 U1718 ( .ip1(n1341), .ip2(n1336), .op(n1339) );
  nand2_1 U1719 ( .ip1(n1337), .ip2(\mult/counterQ [5]), .op(n1338) );
  nand2_1 U1720 ( .ip1(n1339), .ip2(n1338), .op(n631) );
  nand2_1 U1721 ( .ip1(n1341), .ip2(n1797), .op(n1347) );
  inv_1 U1722 ( .ip(n1796), .op(n1787) );
  nor2_1 U1723 ( .ip1(n1787), .ip2(n1342), .op(n1345) );
  nor2_1 U1724 ( .ip1(n1976), .ip2(n1343), .op(n1344) );
  nor2_1 U1725 ( .ip1(n1345), .ip2(n1344), .op(n1346) );
  nand2_1 U1726 ( .ip1(n1347), .ip2(n1346), .op(n629) );
  nand2_1 U1727 ( .ip1(n1293), .ip2(multQ[15]), .op(n1349) );
  nand2_1 U1728 ( .ip1(result2[15]), .ip2(n1354), .op(n1348) );
  nand2_1 U1729 ( .ip1(n1349), .ip2(n1348), .op(n546) );
  nand2_1 U1730 ( .ip1(n1293), .ip2(multQ[14]), .op(n1351) );
  nand2_1 U1731 ( .ip1(result2[14]), .ip2(n1354), .op(n1350) );
  nand2_1 U1732 ( .ip1(n1351), .ip2(n1350), .op(n547) );
  nand2_1 U1733 ( .ip1(n1293), .ip2(multQ[12]), .op(n1353) );
  nand2_1 U1734 ( .ip1(result2[12]), .ip2(n1354), .op(n1352) );
  nand2_1 U1735 ( .ip1(n1353), .ip2(n1352), .op(n549) );
  nand2_1 U1736 ( .ip1(n2064), .ip2(multQ[1]), .op(n1356) );
  nand2_1 U1737 ( .ip1(result2[1]), .ip2(n2049), .op(n1355) );
  nand2_1 U1738 ( .ip1(n1356), .ip2(n1355), .op(n560) );
  nand2_1 U1739 ( .ip1(n1293), .ip2(multQ[10]), .op(n1358) );
  nand2_1 U1740 ( .ip1(result2[10]), .ip2(n1354), .op(n1357) );
  nand2_1 U1741 ( .ip1(n1358), .ip2(n1357), .op(n551) );
  nor2_1 U1742 ( .ip1(partialQ[0]), .ip2(n1359), .op(n1360) );
  nor2_1 U1743 ( .ip1(n2069), .ip2(n1360), .op(n1362) );
  nand2_1 U1744 ( .ip1(n1362), .ip2(n1361), .op(n1364) );
  nand2_1 U1745 ( .ip1(n2064), .ip2(partialQ[0]), .op(n1363) );
  nand2_1 U1746 ( .ip1(n1364), .ip2(n1363), .op(n545) );
  nand2_1 U1747 ( .ip1(n1293), .ip2(multQ[9]), .op(n1366) );
  nand2_1 U1748 ( .ip1(result2[9]), .ip2(n1354), .op(n1365) );
  nand2_1 U1749 ( .ip1(n1366), .ip2(n1365), .op(n552) );
  nand2_1 U1750 ( .ip1(n1293), .ip2(multQ[13]), .op(n1368) );
  nand2_1 U1751 ( .ip1(result2[13]), .ip2(n1354), .op(n1367) );
  nand2_1 U1752 ( .ip1(n1368), .ip2(n1367), .op(n548) );
  nand2_1 U1753 ( .ip1(n1293), .ip2(multQ[11]), .op(n1370) );
  nand2_1 U1754 ( .ip1(result2[11]), .ip2(n1354), .op(n1369) );
  nand2_1 U1755 ( .ip1(n1370), .ip2(n1369), .op(n550) );
  nand2_1 U1756 ( .ip1(n2064), .ip2(multQ[0]), .op(n1372) );
  nand2_1 U1757 ( .ip1(result2[0]), .ip2(n2049), .op(n1371) );
  nand2_1 U1758 ( .ip1(n1372), .ip2(n1371), .op(n561) );
  nand2_1 U1759 ( .ip1(n1293), .ip2(multQ[3]), .op(n1374) );
  nand2_1 U1760 ( .ip1(result2[3]), .ip2(n2059), .op(n1373) );
  nand2_1 U1761 ( .ip1(n1374), .ip2(n1373), .op(n558) );
  nand2_1 U1762 ( .ip1(n1293), .ip2(multQ[7]), .op(n1376) );
  nand2_1 U1763 ( .ip1(result2[7]), .ip2(n2059), .op(n1375) );
  nand2_1 U1764 ( .ip1(n1376), .ip2(n1375), .op(n554) );
  nand2_1 U1765 ( .ip1(n1293), .ip2(multQ[8]), .op(n1378) );
  nand2_1 U1766 ( .ip1(result2[8]), .ip2(n2024), .op(n1377) );
  nand2_1 U1767 ( .ip1(n1378), .ip2(n1377), .op(n553) );
  nand2_1 U1768 ( .ip1(n1293), .ip2(multQ[5]), .op(n1380) );
  nand2_1 U1769 ( .ip1(result2[5]), .ip2(n2059), .op(n1379) );
  nand2_1 U1770 ( .ip1(n1380), .ip2(n1379), .op(n556) );
  nand2_1 U1771 ( .ip1(n1293), .ip2(multQ[4]), .op(n1382) );
  nand2_1 U1772 ( .ip1(result2[4]), .ip2(n2059), .op(n1381) );
  nand2_1 U1773 ( .ip1(n1382), .ip2(n1381), .op(n557) );
  nand2_1 U1774 ( .ip1(n1293), .ip2(multQ[2]), .op(n1384) );
  nand2_1 U1775 ( .ip1(result2[2]), .ip2(n2059), .op(n1383) );
  nand2_1 U1776 ( .ip1(n1384), .ip2(n1383), .op(n559) );
  nand2_1 U1777 ( .ip1(n1293), .ip2(multQ[6]), .op(n1386) );
  nand2_1 U1778 ( .ip1(result2[6]), .ip2(n2059), .op(n1385) );
  nand2_1 U1779 ( .ip1(n1386), .ip2(n1385), .op(n555) );
  nand2_1 U1780 ( .ip1(n1387), .ip2(ramAQ[14]), .op(n1388) );
  nand2_1 U1781 ( .ip1(n1388), .ip2(n2193), .op(n681) );
  nand2_1 U1782 ( .ip1(n1387), .ip2(ramAQ[9]), .op(n1389) );
  nand2_1 U1783 ( .ip1(n1389), .ip2(n2188), .op(n676) );
  nand2_1 U1784 ( .ip1(n1387), .ip2(ramAQ[10]), .op(n1390) );
  nand2_1 U1785 ( .ip1(n1390), .ip2(n2189), .op(n677) );
  nand2_1 U1786 ( .ip1(n1387), .ip2(ramAQ[7]), .op(n1391) );
  nand2_1 U1787 ( .ip1(n1391), .ip2(n2187), .op(n674) );
  nand2_1 U1788 ( .ip1(n1387), .ip2(ramAQ[11]), .op(n1392) );
  nand2_1 U1789 ( .ip1(n1392), .ip2(n2190), .op(n678) );
  nand2_1 U1790 ( .ip1(n1387), .ip2(ramAQ[12]), .op(n1393) );
  nand2_1 U1791 ( .ip1(n1393), .ip2(n2191), .op(n679) );
  nand2_1 U1792 ( .ip1(n1387), .ip2(ramAQ[15]), .op(n1394) );
  nand2_1 U1793 ( .ip1(n1394), .ip2(n2194), .op(n682) );
  nand2_1 U1794 ( .ip1(n1387), .ip2(ramAQ[13]), .op(n1395) );
  nand2_1 U1795 ( .ip1(n1395), .ip2(n2192), .op(n680) );
  inv_1 U1796 ( .ip(counterQ[15]), .op(n1413) );
  inv_1 U1797 ( .ip(counterQ[8]), .op(n2045) );
  inv_1 U1798 ( .ip(n2045), .op(n1444) );
  inv_1 U1799 ( .ip(counterQ[9]), .op(n2048) );
  inv_1 U1800 ( .ip(n2048), .op(n2051) );
  nand2_1 U1801 ( .ip1(n1444), .ip2(n2051), .op(n1452) );
  inv_1 U1802 ( .ip(counterQ[10]), .op(n1449) );
  inv_1 U1803 ( .ip(n1449), .op(n1396) );
  nand2_1 U1804 ( .ip1(n1396), .ip2(counterQ[11]), .op(n1397) );
  nor2_2 U1805 ( .ip1(n1452), .ip2(n1397), .op(n2038) );
  inv_1 U1806 ( .ip(counterQ[12]), .op(n1463) );
  inv_1 U1807 ( .ip(counterQ[13]), .op(n1398) );
  nand2_1 U1808 ( .ip1(n717), .ip2(n2042), .op(n1428) );
  inv_1 U1809 ( .ip(counterQ[14]), .op(n1433) );
  nor2_1 U1810 ( .ip1(n1428), .ip2(n1433), .op(n1399) );
  nand2_1 U1811 ( .ip1(n2038), .ip2(n1399), .op(n1410) );
  inv_1 U1812 ( .ip(counterQ[4]), .op(n1400) );
  inv_1 U1813 ( .ip(counterQ[5]), .op(n1401) );
  nand2_1 U1814 ( .ip1(n1999), .ip2(n1420), .op(n2005) );
  inv_1 U1815 ( .ip(counterQ[6]), .op(n2008) );
  inv_1 U1816 ( .ip(n2008), .op(n1403) );
  inv_1 U1817 ( .ip(counterQ[7]), .op(n1989) );
  inv_1 U1818 ( .ip(n1989), .op(n1402) );
  nand2_1 U1819 ( .ip1(n1403), .ip2(n1402), .op(n1404) );
  nor2_1 U1820 ( .ip1(n2005), .ip2(n1404), .op(n1409) );
  inv_1 U1821 ( .ip(counterQ[3]), .op(n1992) );
  inv_1 U1822 ( .ip(counterQ[2]), .op(n1425) );
  inv_1 U1823 ( .ip(n1425), .op(n1405) );
  nand2_1 U1824 ( .ip1(n1406), .ip2(n1405), .op(n1408) );
  inv_1 U1825 ( .ip(counterQ[1]), .op(n1437) );
  inv_1 U1826 ( .ip(n1437), .op(n1407) );
  nand2_1 U1827 ( .ip1(n1407), .ip2(counterQ[0]), .op(n1423) );
  nand2_2 U1828 ( .ip1(n1409), .ip2(n1417), .op(n2046) );
  nor2_1 U1829 ( .ip1(n1410), .ip2(n2046), .op(n1411) );
  nand2_1 U1830 ( .ip1(n1412), .ip2(n2059), .op(n1416) );
  inv_1 U1831 ( .ip(n1413), .op(n1414) );
  nand2_1 U1832 ( .ip1(n1293), .ip2(n1414), .op(n1415) );
  nand2_1 U1833 ( .ip1(n1416), .ip2(n1415), .op(n635) );
  nor2_1 U1834 ( .ip1(n2006), .ip2(n1400), .op(n1418) );
  nand2_1 U1835 ( .ip1(n1419), .ip2(n2049), .op(n1422) );
  inv_1 U1836 ( .ip(n1401), .op(n1420) );
  nand2_1 U1837 ( .ip1(n2064), .ip2(n1420), .op(n1421) );
  nand2_1 U1838 ( .ip1(n1422), .ip2(n1421), .op(n645) );
  inv_1 U1839 ( .ip(n1423), .op(n1993) );
  nand2_1 U1840 ( .ip1(n1424), .ip2(n2049), .op(n1427) );
  nand2_1 U1841 ( .ip1(n2064), .ip2(n1405), .op(n1426) );
  nand2_1 U1842 ( .ip1(n1427), .ip2(n1426), .op(n648) );
  nand2_1 U1843 ( .ip1(n2038), .ip2(n1429), .op(n1430) );
  nor2_1 U1844 ( .ip1(n1430), .ip2(n2046), .op(n1431) );
  nand2_1 U1845 ( .ip1(n1432), .ip2(n2049), .op(n1436) );
  inv_1 U1846 ( .ip(n1433), .op(n1434) );
  nand2_1 U1847 ( .ip1(n2064), .ip2(n1434), .op(n1435) );
  nand2_1 U1848 ( .ip1(n1436), .ip2(n1435), .op(n636) );
  nand2_1 U1849 ( .ip1(n2064), .ip2(n1407), .op(n1440) );
  nand2_1 U1850 ( .ip1(n1438), .ip2(n2049), .op(n1439) );
  nand2_1 U1851 ( .ip1(n1440), .ip2(n1439), .op(n649) );
  inv_1 U1852 ( .ip(n2208), .op(n1441) );
  nor2_1 U1853 ( .ip1(n1441), .ip2(n2203), .op(n2206) );
  inv_1 U1854 ( .ip(n2224), .op(n1442) );
  nor2_1 U1855 ( .ip1(n1442), .ip2(n2219), .op(n2222) );
  nand2_1 U1856 ( .ip1(n2064), .ip2(n1444), .op(n1445) );
  nand2_1 U1857 ( .ip1(n1446), .ip2(n1445), .op(n642) );
  nor2_1 U1858 ( .ip1(n2046), .ip2(n1452), .op(n1447) );
  nand2_1 U1859 ( .ip1(n1448), .ip2(n1354), .op(n1451) );
  nand2_1 U1860 ( .ip1(n2064), .ip2(n1396), .op(n1450) );
  nand2_1 U1861 ( .ip1(n1451), .ip2(n1450), .op(n640) );
  inv_1 U1862 ( .ip(n1452), .op(n1453) );
  nand2_1 U1863 ( .ip1(n1453), .ip2(n1396), .op(n1454) );
  nor2_1 U1864 ( .ip1(n2046), .ip2(n1454), .op(n1455) );
  nand2_1 U1865 ( .ip1(n1457), .ip2(n1354), .op(n1459) );
  nand2_1 U1866 ( .ip1(n2064), .ip2(counterQ[11]), .op(n1458) );
  nand2_1 U1867 ( .ip1(n1459), .ip2(n1458), .op(n639) );
  inv_1 U1868 ( .ip(n2038), .op(n1460) );
  nor2_1 U1869 ( .ip1(n2046), .ip2(n1460), .op(n1461) );
  nand2_1 U1870 ( .ip1(n1462), .ip2(n2024), .op(n1465) );
  nand2_1 U1871 ( .ip1(n2064), .ip2(n717), .op(n1464) );
  nand2_1 U1872 ( .ip1(n1465), .ip2(n1464), .op(n638) );
  inv_1 U1873 ( .ip(n1487), .op(n1473) );
  inv_1 U1874 ( .ip(n1466), .op(n1472) );
  or2_1 U1875 ( .ip1(n1468), .ip2(n1467), .op(n1469) );
  nor2_2 U1876 ( .ip1(n1472), .ip2(n1471), .op(n1489) );
  nor2_2 U1877 ( .ip1(n1473), .ip2(n1489), .op(n1477) );
  nand2_1 U1878 ( .ip1(n1474), .ip2(n1500), .op(n1475) );
  inv_1 U1879 ( .ip(n1475), .op(n1478) );
  nor2_1 U1880 ( .ip1(n2069), .ip2(n1478), .op(n1476) );
  nand2_1 U1881 ( .ip1(n1477), .ip2(n1476), .op(n1486) );
  inv_1 U1882 ( .ip(n1477), .op(n1480) );
  nor3_1 U1883 ( .ip1(n1481), .ip2(n2069), .ip3(n1475), .op(n1479) );
  nand2_1 U1884 ( .ip1(n1480), .ip2(n1479), .op(n1485) );
  nand2_1 U1885 ( .ip1(n1293), .ip2(partialQ[3]), .op(n1484) );
  inv_1 U1886 ( .ip(n1481), .op(n1488) );
  nor2_1 U1887 ( .ip1(n2069), .ip2(n1488), .op(n1482) );
  nand2_1 U1888 ( .ip1(n1475), .ip2(n1482), .op(n1483) );
  nand4_1 U1889 ( .ip1(n1486), .ip2(n1485), .ip3(n1484), .ip4(n1483), .op(n542) );
  and2_1 U1890 ( .ip1(n1488), .ip2(n1487), .op(n1490) );
  nand2_1 U1891 ( .ip1(n1293), .ip2(partialQ[2]), .op(n1492) );
  nand2_1 U1892 ( .ip1(n1493), .ip2(n1492), .op(n543) );
  inv_1 U1893 ( .ip(n1494), .op(n2076) );
  inv_1 U1894 ( .ip(n1719), .op(n1495) );
  nand2_1 U1895 ( .ip1(n2076), .ip2(n1495), .op(n1497) );
  nand2_1 U1896 ( .ip1(n721), .ip2(\mult/storeQ [0]), .op(n1496) );
  nand2_1 U1897 ( .ip1(n1497), .ip2(n1496), .op(n625) );
  nand2_1 U1898 ( .ip1(n1499), .ip2(n1498), .op(n1503) );
  nand2_2 U1899 ( .ip1(n1501), .ip2(n1500), .op(n1864) );
  inv_2 U1900 ( .ip(n1864), .op(n1502) );
  nand2_4 U1901 ( .ip1(n1502), .ip2(n1503), .op(n2066) );
  buf_1 U1902 ( .ip(n1505), .op(n2058) );
  and2_1 U1903 ( .ip1(n2065), .ip2(n2058), .op(n1506) );
  nand2_1 U1904 ( .ip1(n2066), .ip2(n1506), .op(n1522) );
  buf_1 U1905 ( .ip(n1507), .op(n2056) );
  nor2_1 U1906 ( .ip1(multQ[6]), .ip2(partialQ[6]), .op(n1511) );
  inv_1 U1907 ( .ip(n1508), .op(n2055) );
  nor2_1 U1908 ( .ip1(n1509), .ip2(n2055), .op(n1510) );
  nor2_1 U1909 ( .ip1(n1511), .ip2(n1510), .op(n1512) );
  nor2_1 U1910 ( .ip1(n2056), .ip2(n1512), .op(n1518) );
  nand2_1 U1911 ( .ip1(n1513), .ip2(n1514), .op(n1517) );
  nor2_1 U1912 ( .ip1(n2069), .ip2(n1517), .op(n1515) );
  nand3_1 U1913 ( .ip1(n1522), .ip2(n1518), .ip3(n1515), .op(n1527) );
  nor2_1 U1914 ( .ip1(n1516), .ip2(n1917), .op(n1521) );
  and2_1 U1915 ( .ip1(n1517), .ip2(n2049), .op(n1523) );
  inv_1 U1916 ( .ip(n1523), .op(n1519) );
  nor2_1 U1917 ( .ip1(n1519), .ip2(n1518), .op(n1520) );
  nor2_1 U1918 ( .ip1(n1521), .ip2(n1520), .op(n1526) );
  inv_1 U1919 ( .ip(n1522), .op(n1524) );
  nand2_1 U1920 ( .ip1(n1524), .ip2(n1523), .op(n1525) );
  nand3_1 U1921 ( .ip1(n1527), .ip2(n1526), .ip3(n1525), .op(n538) );
  nand2_2 U1922 ( .ip1(n1529), .ip2(n1528), .op(n1793) );
  or2_1 U1923 ( .ip1(n1530), .ip2(n708), .op(n1534) );
  or2_1 U1924 ( .ip1(n1531), .ip2(n1632), .op(n1533) );
  or2_1 U1925 ( .ip1(n1614), .ip2(n1626), .op(n1532) );
  nand3_2 U1926 ( .ip1(n1534), .ip2(n1533), .ip3(n1532), .op(n1771) );
  inv_2 U1927 ( .ip(n1771), .op(n1686) );
  nor2_1 U1928 ( .ip1(ramAQ[5]), .ip2(n1632), .op(n1536) );
  nor2_1 U1929 ( .ip1(ramAQ[6]), .ip2(n1626), .op(n1535) );
  nor2_2 U1930 ( .ip1(n1536), .ip2(n1535), .op(n1688) );
  and2_1 U1931 ( .ip1(n877), .ip2(n1537), .op(n1539) );
  nor2_1 U1932 ( .ip1(ramAQ[4]), .ip2(n1624), .op(n1538) );
  nor2_2 U1933 ( .ip1(n1539), .ip2(n1538), .op(n1687) );
  nand2_1 U1934 ( .ip1(n1688), .ip2(n1687), .op(n1540) );
  nor2_2 U1935 ( .ip1(n2081), .ip2(n1541), .op(n1739) );
  nand2_1 U1936 ( .ip1(n1793), .ip2(n1739), .op(n1542) );
  nand2_1 U1937 ( .ip1(n1795), .ip2(n1542), .op(n1560) );
  nor2_1 U1938 ( .ip1(ramAQ[13]), .ip2(n1632), .op(n1544) );
  nor2_1 U1939 ( .ip1(ramAQ[14]), .ip2(n1626), .op(n1543) );
  nor2_1 U1940 ( .ip1(ramAQ[12]), .ip2(n1624), .op(n1546) );
  nor2_1 U1941 ( .ip1(ramAQ[11]), .ip2(n1630), .op(n1545) );
  nand2_1 U1942 ( .ip1(n1770), .ip2(n1796), .op(n1558) );
  nor2_1 U1943 ( .ip1(ramAQ[9]), .ip2(n1632), .op(n1550) );
  nor2_1 U1944 ( .ip1(ramAQ[10]), .ip2(n1626), .op(n1549) );
  nor2_1 U1945 ( .ip1(ramAQ[7]), .ip2(n1630), .op(n1552) );
  nor2_1 U1946 ( .ip1(ramAQ[8]), .ip2(n708), .op(n1551) );
  nand2_1 U1947 ( .ip1(n1772), .ip2(n1978), .op(n1557) );
  nor2_1 U1948 ( .ip1(n1555), .ip2(n1630), .op(n1577) );
  nand2_1 U1949 ( .ip1(n1577), .ip2(n1797), .op(n1556) );
  nand4_1 U1950 ( .ip1(n1802), .ip2(n1558), .ip3(n1557), .ip4(n1556), .op(
        n1559) );
  nand2_1 U1951 ( .ip1(n1560), .ip2(n1559), .op(n1562) );
  nand2_1 U1952 ( .ip1(n1805), .ip2(\mult/storeQ [22]), .op(n1561) );
  nand2_1 U1953 ( .ip1(n1562), .ip2(n1561), .op(n603) );
  nand2_1 U1954 ( .ip1(n1564), .ip2(n1795), .op(n1572) );
  nand2_1 U1955 ( .ip1(n1565), .ip2(n1796), .op(n1570) );
  inv_1 U1956 ( .ip(n1566), .op(n1567) );
  nand2_1 U1957 ( .ip1(n1567), .ip2(n1797), .op(n1569) );
  nand2_1 U1958 ( .ip1(n1722), .ip2(n1978), .op(n1568) );
  nand4_1 U1959 ( .ip1(n1570), .ip2(n1802), .ip3(n1569), .ip4(n1568), .op(
        n1571) );
  nand2_1 U1960 ( .ip1(n2078), .ip2(\mult/storeQ [20]), .op(n1573) );
  nand2_1 U1961 ( .ip1(n1576), .ip2(n1575), .op(n1645) );
  nand2_1 U1962 ( .ip1(n1578), .ip2(n1976), .op(n1581) );
  nand2_1 U1963 ( .ip1(n1688), .ip2(n1687), .op(n1774) );
  nor2_1 U1964 ( .ip1(n1785), .ip2(n1774), .op(n1579) );
  not_ab_or_c_or_d U1965 ( .ip1(n1796), .ip2(n1772), .ip3(\mult/counterQ [4]), 
        .ip4(n1579), .op(n1580) );
  nand2_1 U1966 ( .ip1(n1581), .ip2(n1580), .op(n1583) );
  nand2_1 U1967 ( .ip1(n1686), .ip2(\mult/counterQ [4]), .op(n1582) );
  nand2_1 U1968 ( .ip1(n1583), .ip2(n1582), .op(n1584) );
  inv_1 U1969 ( .ip(n1584), .op(n1585) );
  nand2_1 U1970 ( .ip1(n1645), .ip2(n1585), .op(n1587) );
  nand2_1 U1971 ( .ip1(n2093), .ip2(\mult/storeQ [18]), .op(n1586) );
  nand2_1 U1972 ( .ip1(n1587), .ip2(n1586), .op(n2229) );
  nand2_1 U1973 ( .ip1(n2074), .ip2(\mult/counterQ [4]), .op(n1594) );
  inv_1 U1974 ( .ip(n1786), .op(n1588) );
  nand2_1 U1975 ( .ip1(n1588), .ip2(n1978), .op(n1592) );
  nand2_1 U1976 ( .ip1(n1589), .ip2(n1796), .op(n1591) );
  nand2_1 U1977 ( .ip1(n1783), .ip2(n1797), .op(n1590) );
  nand4_1 U1978 ( .ip1(n1802), .ip2(n1592), .ip3(n1591), .ip4(n1590), .op(
        n1593) );
  and2_1 U1979 ( .ip1(n1594), .ip2(n1593), .op(n1595) );
  nand2_1 U1980 ( .ip1(n1645), .ip2(n1595), .op(n1597) );
  nand2_1 U1981 ( .ip1(n721), .ip2(\mult/storeQ [19]), .op(n1596) );
  nand2_1 U1982 ( .ip1(n1597), .ip2(n1596), .op(n2230) );
  nand2_1 U1983 ( .ip1(n1618), .ip2(ramAQ[1]), .op(n1599) );
  nand2_1 U1984 ( .ip1(n1619), .ip2(ramAQ[0]), .op(n1598) );
  nor2_1 U1985 ( .ip1(n1802), .ip2(n2002), .op(n1643) );
  nand2_1 U1986 ( .ip1(n1613), .ip2(ramAQ[15]), .op(n1602) );
  nand2_1 U1987 ( .ip1(n824), .ip2(ramAQ[14]), .op(n1601) );
  inv_1 U1988 ( .ip(ramAQ[11]), .op(n1603) );
  nor2_1 U1989 ( .ip1(n1603), .ip2(n708), .op(n1606) );
  nor2_1 U1990 ( .ip1(n1604), .ip2(n1626), .op(n1605) );
  inv_1 U1991 ( .ip(ramAQ[10]), .op(n1607) );
  nor2_1 U1992 ( .ip1(n1608), .ip2(n1632), .op(n1609) );
  nand2_1 U1993 ( .ip1(n1613), .ip2(ramAQ[3]), .op(n1617) );
  inv_1 U1994 ( .ip(n1614), .op(n1615) );
  nand2_1 U1995 ( .ip1(n877), .ip2(n1615), .op(n1616) );
  nand2_1 U1996 ( .ip1(n1618), .ip2(ramAQ[5]), .op(n1621) );
  nand2_1 U1997 ( .ip1(n1619), .ip2(ramAQ[4]), .op(n1620) );
  nor2_2 U1998 ( .ip1(n1623), .ip2(n1622), .op(n1975) );
  nor2_1 U1999 ( .ip1(n1785), .ip2(n1975), .op(n1640) );
  inv_1 U2000 ( .ip(ramAQ[7]), .op(n1625) );
  nor2_1 U2001 ( .ip1(n1625), .ip2(n708), .op(n1629) );
  nor2_1 U2002 ( .ip1(n1627), .ip2(n1626), .op(n1628) );
  inv_1 U2003 ( .ip(ramAQ[6]), .op(n1631) );
  nor2_1 U2004 ( .ip1(n1631), .ip2(n1630), .op(n1635) );
  nor2_1 U2005 ( .ip1(n1633), .ip2(n1632), .op(n1634) );
  nand2_1 U2006 ( .ip1(n2083), .ip2(n1796), .op(n1638) );
  nand2_1 U2007 ( .ip1(n1638), .ip2(n1802), .op(n1639) );
  not_ab_or_c_or_d U2008 ( .ip1(n1976), .ip2(n1641), .ip3(n1640), .ip4(n1639), 
        .op(n1642) );
  nor2_1 U2009 ( .ip1(n1643), .ip2(n1642), .op(n1644) );
  nand2_1 U2010 ( .ip1(n1645), .ip2(n1644), .op(n1647) );
  nand2_1 U2011 ( .ip1(n2078), .ip2(\mult/storeQ [17]), .op(n1646) );
  nand2_1 U2012 ( .ip1(n1647), .ip2(n1646), .op(n2231) );
  nand2_1 U2013 ( .ip1(n1832), .ip2(\mult/productQ [11]), .op(n1668) );
  nand2_1 U2014 ( .ip1(n1648), .ip2(n1965), .op(n1661) );
  and2_1 U2015 ( .ip1(n1657), .ip2(n1656), .op(n1966) );
  inv_1 U2016 ( .ip(n1966), .op(n1658) );
  nor3_1 U2017 ( .ip1(n1659), .ip2(n1660), .ip3(n1658), .op(n1664) );
  nand3_1 U2018 ( .ip1(n1661), .ip2(n1964), .ip3(n1660), .op(n1662) );
  nor2_1 U2019 ( .ip1(n1662), .ip2(n1966), .op(n1663) );
  nor3_1 U2020 ( .ip1(n1665), .ip2(n1664), .ip3(n1663), .op(n1666) );
  nand2_1 U2021 ( .ip1(n1666), .ip2(n1856), .op(n1667) );
  nand2_1 U2022 ( .ip1(n1668), .ip2(n1667), .op(n582) );
  and2_1 U2023 ( .ip1(n1786), .ip2(\mult/counterQ [2]), .op(n1673) );
  nand2_1 U2024 ( .ip1(n1669), .ip2(n1973), .op(n1671) );
  nand2_1 U2025 ( .ip1(n2074), .ip2(n2081), .op(n1670) );
  nand2_1 U2026 ( .ip1(n1671), .ip2(n1670), .op(n1672) );
  nand2_1 U2027 ( .ip1(n1675), .ip2(n1674), .op(n1676) );
  nand2_1 U2028 ( .ip1(n1677), .ip2(n1676), .op(n614) );
  nand2_1 U2029 ( .ip1(n1730), .ip2(n2081), .op(n1682) );
  and2_1 U2030 ( .ip1(n1678), .ip2(n1973), .op(n1680) );
  nor2_1 U2031 ( .ip1(n2084), .ip2(n1722), .op(n1679) );
  and2_1 U2032 ( .ip1(n1682), .ip2(n1681), .op(n1683) );
  nand2_1 U2033 ( .ip1(n2092), .ip2(n1683), .op(n1685) );
  nand2_1 U2034 ( .ip1(n1805), .ip2(\mult/storeQ [12]), .op(n1684) );
  nand2_1 U2035 ( .ip1(n1685), .ip2(n1684), .op(n613) );
  and2_1 U2036 ( .ip1(n1686), .ip2(n2081), .op(n1693) );
  nor2_1 U2037 ( .ip1(n2086), .ip2(n1772), .op(n1692) );
  nand2_1 U2038 ( .ip1(n1688), .ip2(n1687), .op(n1689) );
  nand2_1 U2039 ( .ip1(n1689), .ip2(\mult/counterQ [2]), .op(n1690) );
  nand2_1 U2040 ( .ip1(n1690), .ip2(n1785), .op(n1691) );
  nand2_1 U2041 ( .ip1(n2092), .ip2(n1694), .op(n1696) );
  nand2_1 U2042 ( .ip1(n2078), .ip2(\mult/storeQ [10]), .op(n1695) );
  nand2_1 U2043 ( .ip1(n1696), .ip2(n1695), .op(n615) );
  nand2_1 U2044 ( .ip1(n1702), .ip2(n1701), .op(n1697) );
  nand2_1 U2045 ( .ip1(n1697), .ip2(n1354), .op(n1698) );
  inv_1 U2046 ( .ip(n1698), .op(n1714) );
  buf_1 U2047 ( .ip(n1699), .op(n1711) );
  inv_1 U2048 ( .ip(n1711), .op(n1708) );
  nor2_1 U2049 ( .ip1(n1700), .ip2(n1917), .op(n1707) );
  nor2_2 U2050 ( .ip1(n1704), .ip2(n1703), .op(n1902) );
  nor2_1 U2051 ( .ip1(n1902), .ip2(n1705), .op(n1706) );
  not_ab_or_c_or_d U2052 ( .ip1(n1714), .ip2(n1708), .ip3(n1707), .ip4(n1706), 
        .op(n1718) );
  buf_1 U2053 ( .ip(n1709), .op(n1713) );
  nor2_1 U2054 ( .ip1(n2069), .ip2(n1710), .op(n1712) );
  nand4_1 U2055 ( .ip1(n1713), .ip2(n1902), .ip3(n1712), .ip4(n1711), .op(
        n1717) );
  inv_1 U2056 ( .ip(n1713), .op(n1715) );
  nand2_1 U2057 ( .ip1(n1715), .ip2(n1714), .op(n1716) );
  nand3_1 U2058 ( .ip1(n1718), .ip2(n1717), .ip3(n1716), .op(n537) );
  nand2_1 U2059 ( .ip1(n1719), .ip2(n2081), .op(n1720) );
  nand2_1 U2060 ( .ip1(n1720), .ip2(n1785), .op(n1725) );
  and2_1 U2061 ( .ip1(\mult/counterQ [2]), .ip2(n1721), .op(n1724) );
  nor2_1 U2062 ( .ip1(n2086), .ip2(n1722), .op(n1723) );
  nand2_1 U2063 ( .ip1(n2092), .ip2(n1726), .op(n1729) );
  nand2_1 U2064 ( .ip1(n721), .ip2(\mult/storeQ [8]), .op(n1728) );
  nand2_1 U2065 ( .ip1(n1729), .ip2(n1728), .op(n617) );
  nor2_1 U2066 ( .ip1(n2081), .ip2(n1730), .op(n1731) );
  nand2_1 U2067 ( .ip1(n2092), .ip2(n1731), .op(n1733) );
  nand2_1 U2068 ( .ip1(n721), .ip2(\mult/storeQ [4]), .op(n1732) );
  nand2_1 U2069 ( .ip1(n1733), .ip2(n1732), .op(n621) );
  inv_1 U2070 ( .ip(n2002), .op(n1735) );
  nand2_1 U2071 ( .ip1(n2092), .ip2(n1792), .op(n1738) );
  nand2_1 U2072 ( .ip1(n1805), .ip2(\mult/storeQ [5]), .op(n1737) );
  nand2_1 U2073 ( .ip1(n1738), .ip2(n1737), .op(n620) );
  nand2_1 U2074 ( .ip1(n2092), .ip2(n1739), .op(n1741) );
  nand2_1 U2075 ( .ip1(n1727), .ip2(\mult/storeQ [6]), .op(n1740) );
  nand2_1 U2076 ( .ip1(n1741), .ip2(n1740), .op(n619) );
  nand2_1 U2077 ( .ip1(n1743), .ip2(n1742), .op(n1744) );
  and2_1 U2078 ( .ip1(n2066), .ip2(n1744), .op(n1754) );
  inv_1 U2079 ( .ip(n1745), .op(n1746) );
  and2_1 U2080 ( .ip1(n713), .ip2(n1749), .op(n1747) );
  nor2_2 U2081 ( .ip1(n1747), .ip2(n2054), .op(n1755) );
  nor2_1 U2082 ( .ip1(n2069), .ip2(n1755), .op(n1748) );
  nand2_1 U2083 ( .ip1(n1754), .ip2(n1748), .op(n1762) );
  nor2_1 U2084 ( .ip1(n1749), .ip2(n1917), .op(n1753) );
  inv_1 U2085 ( .ip(n1750), .op(n1751) );
  nand2_1 U2086 ( .ip1(n1125), .ip2(n1751), .op(n1763) );
  nor3_1 U2087 ( .ip1(n1763), .ip2(n2069), .ip3(n1755), .op(n1752) );
  nor2_1 U2088 ( .ip1(n1753), .ip2(n1752), .op(n1761) );
  inv_1 U2089 ( .ip(n1754), .op(n1759) );
  nand2_1 U2090 ( .ip1(n1763), .ip2(n2059), .op(n1757) );
  inv_1 U2091 ( .ip(n1755), .op(n1756) );
  nand2_1 U2092 ( .ip1(n1759), .ip2(n1758), .op(n1760) );
  nand3_1 U2093 ( .ip1(n1762), .ip2(n1761), .ip3(n1760), .op(n540) );
  and2_1 U2094 ( .ip1(n1763), .ip2(n1744), .op(n1764) );
  xor2_1 U2095 ( .ip1(n1764), .ip2(n2066), .op(n1765) );
  nand2_4 U2096 ( .ip1(n1765), .ip2(n2059), .op(n1767) );
  nand2_1 U2097 ( .ip1(n1293), .ip2(partialQ[4]), .op(n1766) );
  nand2_1 U2098 ( .ip1(n1767), .ip2(n1766), .op(n541) );
  nand2_1 U2099 ( .ip1(n2076), .ip2(n1771), .op(n1769) );
  nand2_1 U2100 ( .ip1(n721), .ip2(\mult/storeQ [2]), .op(n1768) );
  nand2_1 U2101 ( .ip1(n1769), .ip2(n1768), .op(n623) );
  nor2_1 U2102 ( .ip1(n2086), .ip2(n1770), .op(n1779) );
  nor2_1 U2103 ( .ip1(n1785), .ip2(n1771), .op(n1778) );
  nand2_1 U2104 ( .ip1(n1773), .ip2(n1797), .op(n1776) );
  nand2_1 U2105 ( .ip1(n1774), .ip2(n1796), .op(n1775) );
  nand2_1 U2106 ( .ip1(n2092), .ip2(n1780), .op(n1782) );
  nand2_1 U2107 ( .ip1(n1805), .ip2(\mult/storeQ [14]), .op(n1781) );
  nand2_1 U2108 ( .ip1(n1782), .ip2(n1781), .op(n611) );
  nand2_1 U2109 ( .ip1(n1783), .ip2(n1976), .op(n1784) );
  nand2_1 U2110 ( .ip1(n1784), .ip2(n2084), .op(n1791) );
  nor2_1 U2111 ( .ip1(n1785), .ip2(n2074), .op(n1789) );
  nor2_1 U2112 ( .ip1(n1787), .ip2(n1786), .op(n1788) );
  nand2_1 U2113 ( .ip1(n1793), .ip2(n1792), .op(n1794) );
  nand2_1 U2114 ( .ip1(n1795), .ip2(n1794), .op(n1804) );
  nand2_1 U2115 ( .ip1(n2085), .ip2(n1796), .op(n1801) );
  nand2_1 U2116 ( .ip1(n2083), .ip2(n1978), .op(n1800) );
  nand2_1 U2117 ( .ip1(n1798), .ip2(n1797), .op(n1799) );
  nand4_1 U2118 ( .ip1(n1802), .ip2(n1801), .ip3(n1800), .ip4(n1799), .op(
        n1803) );
  nand2_1 U2119 ( .ip1(n1804), .ip2(n1803), .op(n1807) );
  nand2_1 U2120 ( .ip1(n1805), .ip2(\mult/storeQ [21]), .op(n1806) );
  nand2_1 U2121 ( .ip1(n1807), .ip2(n1806), .op(n604) );
  nand2_1 U2122 ( .ip1(n1808), .ip2(\mult/productQ [12]), .op(n1818) );
  or2_1 U2123 ( .ip1(n1810), .ip2(n1809), .op(n1815) );
  nand2_1 U2124 ( .ip1(n1812), .ip2(n1811), .op(n1942) );
  inv_1 U2125 ( .ip(n1942), .op(n1813) );
  nand2_1 U2126 ( .ip1(n1954), .ip2(n1813), .op(n1814) );
  xnor2_1 U2127 ( .ip1(n1815), .ip2(n1814), .op(n1816) );
  nand2_1 U2128 ( .ip1(n1816), .ip2(n1856), .op(n1817) );
  nand2_1 U2129 ( .ip1(n1818), .ip2(n1817), .op(n581) );
  nor2_1 U2130 ( .ip1(\mult/storeQ [20]), .ip2(\mult/productQ [20]), .op(n1844) );
  inv_1 U2131 ( .ip(n1844), .op(n2144) );
  nand2_1 U2132 ( .ip1(\mult/productQ [20]), .ip2(\mult/storeQ [20]), .op(
        n2142) );
  and2_1 U2133 ( .ip1(n2144), .ip2(n2142), .op(n1828) );
  or2_1 U2134 ( .ip1(\mult/storeQ [17]), .ip2(\mult/productQ [17]), .op(n2097)
         );
  nand2_1 U2135 ( .ip1(n2097), .ip2(n2101), .op(n1819) );
  nand2_1 U2136 ( .ip1(\mult/storeQ [17]), .ip2(\mult/productQ [17]), .op(
        n2096) );
  or2_1 U2137 ( .ip1(\mult/storeQ [18]), .ip2(\mult/productQ [18]), .op(n2113)
         );
  or2_1 U2138 ( .ip1(\mult/storeQ [19]), .ip2(\mult/productQ [19]), .op(n2108)
         );
  nand2_1 U2139 ( .ip1(n2113), .ip2(n2108), .op(n1825) );
  inv_1 U2140 ( .ip(n1825), .op(n1820) );
  nand2_1 U2141 ( .ip1(n2110), .ip2(n1820), .op(n1824) );
  and2_1 U2142 ( .ip1(\mult/productQ [19]), .ip2(\mult/storeQ [19]), .op(n2107) );
  nand2_1 U2143 ( .ip1(\mult/storeQ [18]), .ip2(\mult/productQ [18]), .op(
        n2111) );
  inv_1 U2144 ( .ip(n2108), .op(n1821) );
  nor2_1 U2145 ( .ip1(n2111), .ip2(n1821), .op(n1822) );
  nor2_1 U2146 ( .ip1(n2107), .ip2(n1822), .op(n1823) );
  nand2_1 U2147 ( .ip1(n2098), .ip2(n2097), .op(n2115) );
  inv_1 U2148 ( .ip(n2145), .op(n1851) );
  nor2_1 U2149 ( .ip1(n1851), .ip2(n2126), .op(n1826) );
  nor2_1 U2150 ( .ip1(n2141), .ip2(n1826), .op(n1827) );
  nand2_1 U2151 ( .ip1(n1829), .ip2(n1856), .op(n1831) );
  nand2_1 U2152 ( .ip1(n2123), .ip2(\mult/productQ [20]), .op(n1830) );
  nand2_1 U2153 ( .ip1(n1831), .ip2(n1830), .op(n573) );
  nand2_1 U2154 ( .ip1(n1832), .ip2(\mult/productQ [18]), .op(n1840) );
  and2_1 U2155 ( .ip1(n2113), .ip2(n2111), .op(n1837) );
  nor2_2 U2156 ( .ip1(n1834), .ip2(n1833), .op(n2146) );
  nor2_1 U2157 ( .ip1(n2146), .ip2(n2115), .op(n1835) );
  nor2_1 U2158 ( .ip1(n2110), .ip2(n1835), .op(n1836) );
  xnor2_1 U2159 ( .ip1(n1837), .ip2(n1836), .op(n1838) );
  nand2_1 U2160 ( .ip1(n1838), .ip2(n1856), .op(n1839) );
  nand2_1 U2161 ( .ip1(n1840), .ip2(n1839), .op(n575) );
  nand2_1 U2162 ( .ip1(n1841), .ip2(\mult/productQ [23]), .op(n1859) );
  nand2_1 U2163 ( .ip1(\mult/productQ [23]), .ip2(\mult/storeQ [23]), .op(
        n1843) );
  or2_1 U2164 ( .ip1(\mult/storeQ [23]), .ip2(\mult/productQ [23]), .op(n1842)
         );
  and2_1 U2165 ( .ip1(n1843), .ip2(n1842), .op(n1855) );
  nor2_1 U2166 ( .ip1(\mult/storeQ [21]), .ip2(\mult/productQ [21]), .op(n2139) );
  nor2_1 U2167 ( .ip1(n1844), .ip2(n2139), .op(n2128) );
  or2_1 U2168 ( .ip1(\mult/storeQ [22]), .ip2(\mult/productQ [22]), .op(n2125)
         );
  nand2_1 U2169 ( .ip1(n2128), .ip2(n2125), .op(n1850) );
  nand2_1 U2170 ( .ip1(n2141), .ip2(n1845), .op(n1849) );
  nand2_1 U2171 ( .ip1(\mult/productQ [22]), .ip2(\mult/storeQ [22]), .op(
        n2124) );
  and2_1 U2172 ( .ip1(\mult/productQ [21]), .ip2(\mult/storeQ [21]), .op(n2138) );
  nor2_1 U2173 ( .ip1(n2142), .ip2(n2139), .op(n1846) );
  nand2_1 U2174 ( .ip1(n1847), .ip2(n2125), .op(n1848) );
  nand3_1 U2175 ( .ip1(n1849), .ip2(n2124), .ip3(n1848), .op(n1853) );
  nor2_1 U2176 ( .ip1(n2146), .ip2(n744), .op(n1852) );
  nor2_1 U2177 ( .ip1(n1853), .ip2(n1852), .op(n1854) );
  nand2_1 U2178 ( .ip1(n1859), .ip2(n1858), .op(n570) );
  nand2_1 U2179 ( .ip1(n2012), .ip2(n1899), .op(n1860) );
  inv_1 U2180 ( .ip(n1860), .op(n1869) );
  nor2_1 U2181 ( .ip1(n1861), .ip2(n1862), .op(n1868) );
  nand2_1 U2182 ( .ip1(n1864), .ip2(n1863), .op(n1903) );
  or2_1 U2183 ( .ip1(n1866), .ip2(n1865), .op(n1867) );
  nand3_1 U2184 ( .ip1(n1868), .ip2(n1903), .ip3(n1867), .op(n1927) );
  nand2_1 U2185 ( .ip1(n1869), .ip2(n1927), .op(n1893) );
  or2_1 U2186 ( .ip1(n1893), .ip2(n1870), .op(n1896) );
  nand2_1 U2187 ( .ip1(n1872), .ip2(n1871), .op(n1874) );
  nand2_1 U2188 ( .ip1(n1874), .ip2(n1873), .op(n1875) );
  inv_1 U2189 ( .ip(n1875), .op(n2019) );
  or2_1 U2190 ( .ip1(n1877), .ip2(n1876), .op(n2018) );
  nand2_1 U2191 ( .ip1(n2019), .ip2(n2018), .op(n1878) );
  nand2_1 U2192 ( .ip1(n1899), .ip2(n1878), .op(n1879) );
  nand2_1 U2193 ( .ip1(n1879), .ip2(n2016), .op(n1880) );
  nand2_1 U2194 ( .ip1(n1881), .ip2(n1880), .op(n1884) );
  or2_1 U2195 ( .ip1(n1882), .ip2(n1917), .op(n1883) );
  nand2_1 U2196 ( .ip1(n1884), .ip2(n1883), .op(n1885) );
  inv_1 U2197 ( .ip(n1885), .op(n1895) );
  nand2_1 U2198 ( .ip1(n1898), .ip2(n1897), .op(n1886) );
  nand2_1 U2199 ( .ip1(n1899), .ip2(n1886), .op(n1887) );
  nand2_1 U2200 ( .ip1(n1887), .ip2(n2016), .op(n1891) );
  inv_1 U2201 ( .ip(n1888), .op(n1889) );
  or2_1 U2202 ( .ip1(n2069), .ip2(n1889), .op(n1890) );
  nor2_1 U2203 ( .ip1(n1891), .ip2(n1890), .op(n1892) );
  nand2_1 U2204 ( .ip1(n1893), .ip2(n1892), .op(n1894) );
  nand3_1 U2205 ( .ip1(n1895), .ip2(n1896), .ip3(n1894), .op(n532) );
  nand2_1 U2206 ( .ip1(n1898), .ip2(n1897), .op(n1909) );
  nand2_1 U2207 ( .ip1(n2016), .ip2(n1899), .op(n1908) );
  and2_1 U2208 ( .ip1(n1908), .ip2(n2024), .op(n1911) );
  nand2_1 U2209 ( .ip1(n1909), .ip2(n1911), .op(n1901) );
  nand2_1 U2210 ( .ip1(n1293), .ip2(partialQ[12]), .op(n1900) );
  and2_1 U2211 ( .ip1(n1901), .ip2(n1900), .op(n1916) );
  inv_1 U2212 ( .ip(n1905), .op(n1906) );
  nor2_1 U2213 ( .ip1(n1909), .ip2(n743), .op(n1910) );
  nand2_1 U2214 ( .ip1(n1913), .ip2(n1910), .op(n1915) );
  inv_1 U2215 ( .ip(n1911), .op(n1912) );
  or2_1 U2216 ( .ip1(n1913), .ip2(n1912), .op(n1914) );
  nand3_1 U2217 ( .ip1(n1916), .ip2(n1915), .ip3(n1914), .op(n533) );
  nor2_1 U2218 ( .ip1(n1918), .ip2(n1917), .op(n1925) );
  nand2_1 U2219 ( .ip1(n1920), .ip2(n1919), .op(n1933) );
  inv_1 U2220 ( .ip(n1933), .op(n1923) );
  nor2_2 U2221 ( .ip1(n1922), .ip2(n1921), .op(n1931) );
  or2_1 U2222 ( .ip1(n2069), .ip2(n1931), .op(n1926) );
  nor2_1 U2223 ( .ip1(n1926), .ip2(n1923), .op(n1924) );
  nor2_1 U2224 ( .ip1(n1925), .ip2(n1924), .op(n1939) );
  or2_1 U2225 ( .ip1(n1929), .ip2(n1926), .op(n1928) );
  inv_1 U2226 ( .ip(n1927), .op(n1930) );
  or2_1 U2227 ( .ip1(n1928), .ip2(n1930), .op(n1938) );
  or2_1 U2228 ( .ip1(n1930), .ip2(n1929), .op(n1936) );
  inv_1 U2229 ( .ip(n1931), .op(n1932) );
  or3_1 U2230 ( .ip1(n2069), .ip2(n1933), .ip3(n1932), .op(n1934) );
  inv_1 U2231 ( .ip(n1934), .op(n1935) );
  nand2_1 U2232 ( .ip1(n1936), .ip2(n1935), .op(n1937) );
  nand3_1 U2233 ( .ip1(n1938), .ip2(n1939), .ip3(n1937), .op(n535) );
  nand2_1 U2234 ( .ip1(n1808), .ip2(\mult/productQ [14]), .op(n1963) );
  nor2_2 U2235 ( .ip1(n1941), .ip2(n1940), .op(n1955) );
  inv_1 U2236 ( .ip(n1945), .op(n1943) );
  and2_1 U2237 ( .ip1(n1942), .ip2(n1956), .op(n1947) );
  nand2_1 U2238 ( .ip1(n1944), .ip2(n1954), .op(n1953) );
  nor2_1 U2239 ( .ip1(n1956), .ip2(n1955), .op(n1946) );
  mux2_4 U2240 ( .ip1(n1955), .ip2(n1946), .s(n1945), .op(n1951) );
  and2_1 U2241 ( .ip1(n1953), .ip2(n1952), .op(n1959) );
  inv_1 U2242 ( .ip(n1954), .op(n1957) );
  nand3_1 U2243 ( .ip1(n1957), .ip2(n1956), .ip3(n1955), .op(n1958) );
  nand2_1 U2244 ( .ip1(n1959), .ip2(n1958), .op(n1961) );
  or2_1 U2245 ( .ip1(n1961), .ip2(n1960), .op(n1962) );
  nand2_1 U2246 ( .ip1(n1963), .ip2(n1962), .op(n579) );
  nand2_1 U2247 ( .ip1(n2123), .ip2(\mult/productQ [10]), .op(n1972) );
  nand2_1 U2248 ( .ip1(n1965), .ip2(n1964), .op(n1968) );
  nand2_1 U2249 ( .ip1(n1856), .ip2(n1970), .op(n1971) );
  nand2_1 U2250 ( .ip1(n1972), .ip2(n1971), .op(n583) );
  nand2_1 U2251 ( .ip1(n1974), .ip2(n1973), .op(n1981) );
  nand2_1 U2252 ( .ip1(n1975), .ip2(\mult/counterQ [2]), .op(n1980) );
  nor2_1 U2253 ( .ip1(n1976), .ip2(n2002), .op(n1977) );
  nor2_1 U2254 ( .ip1(n1978), .ip2(n1977), .op(n1979) );
  and3_1 U2255 ( .ip1(n1981), .ip2(n1980), .ip3(n1979), .op(n1982) );
  nand2_1 U2256 ( .ip1(n2092), .ip2(n1982), .op(n1984) );
  nand2_1 U2257 ( .ip1(n1727), .ip2(\mult/storeQ [9]), .op(n1983) );
  nand2_1 U2258 ( .ip1(n1984), .ip2(n1983), .op(n616) );
  inv_1 U2259 ( .ip(n2005), .op(n1985) );
  nand2_1 U2260 ( .ip1(n1985), .ip2(n1403), .op(n1986) );
  nand2_1 U2261 ( .ip1(n1988), .ip2(n2049), .op(n1991) );
  nand2_1 U2262 ( .ip1(n2064), .ip2(n1402), .op(n1990) );
  nand2_1 U2263 ( .ip1(n1991), .ip2(n1990), .op(n643) );
  and2_1 U2264 ( .ip1(n1993), .ip2(n1405), .op(n1994) );
  nand2_1 U2265 ( .ip1(n1996), .ip2(n2049), .op(n1998) );
  nand2_1 U2266 ( .ip1(n2064), .ip2(n1406), .op(n1997) );
  nand2_1 U2267 ( .ip1(n1998), .ip2(n1997), .op(n647) );
  inv_1 U2268 ( .ip(n1400), .op(n1999) );
  nand2_1 U2269 ( .ip1(n1999), .ip2(n2064), .op(n2000) );
  nand2_1 U2270 ( .ip1(n2001), .ip2(n2000), .op(n646) );
  nand2_1 U2271 ( .ip1(n2076), .ip2(n2002), .op(n2004) );
  inv_1 U2272 ( .ip(n2077), .op(n2093) );
  nand2_1 U2273 ( .ip1(n2093), .ip2(\mult/storeQ [1]), .op(n2003) );
  nand2_1 U2274 ( .ip1(n2004), .ip2(n2003), .op(n624) );
  nor2_1 U2275 ( .ip1(n2006), .ip2(n2005), .op(n2007) );
  nand2_1 U2276 ( .ip1(n2009), .ip2(n2049), .op(n2011) );
  nand2_1 U2277 ( .ip1(n2064), .ip2(n1403), .op(n2010) );
  nand2_1 U2278 ( .ip1(n2011), .ip2(n2010), .op(n644) );
  and2_1 U2279 ( .ip1(n2012), .ip2(n2020), .op(n2014) );
  nand2_1 U2280 ( .ip1(n2014), .ip2(n2013), .op(n2034) );
  nor2_1 U2281 ( .ip1(n2017), .ip2(n1153), .op(n2029) );
  nand2_1 U2282 ( .ip1(n2019), .ip2(n2018), .op(n2021) );
  nand2_1 U2283 ( .ip1(n2021), .ip2(n2020), .op(n2030) );
  nand2_1 U2284 ( .ip1(n2029), .ip2(n2030), .op(n2026) );
  nand2_1 U2285 ( .ip1(n2023), .ip2(n2022), .op(n2028) );
  nand2_1 U2286 ( .ip1(n2034), .ip2(n2027), .op(n2037) );
  nand2_1 U2287 ( .ip1(n1293), .ip2(partialQ[14]), .op(n2031) );
  nand3_1 U2288 ( .ip1(n2031), .ip2(n2030), .ip3(n2029), .op(n2032) );
  nand2_1 U2289 ( .ip1(n2033), .ip2(n2032), .op(n2036) );
  or2_1 U2290 ( .ip1(n2034), .ip2(n740), .op(n2035) );
  nand3_1 U2291 ( .ip1(n2035), .ip2(n2036), .ip3(n2037), .op(n531) );
  nand2_1 U2292 ( .ip1(n2038), .ip2(n717), .op(n2039) );
  nor2_1 U2293 ( .ip1(n2039), .ip2(n2046), .op(n2040) );
  nand2_1 U2294 ( .ip1(n2041), .ip2(n2049), .op(n2044) );
  inv_1 U2295 ( .ip(n1398), .op(n2042) );
  nand2_1 U2296 ( .ip1(n2064), .ip2(n2042), .op(n2043) );
  nand2_1 U2297 ( .ip1(n2044), .ip2(n2043), .op(n637) );
  nor2_1 U2298 ( .ip1(n2046), .ip2(n2045), .op(n2047) );
  nand2_1 U2299 ( .ip1(n2050), .ip2(n2049), .op(n2053) );
  nand2_1 U2300 ( .ip1(n2064), .ip2(n2051), .op(n2052) );
  nand2_1 U2301 ( .ip1(n2053), .ip2(n2052), .op(n641) );
  or2_1 U2302 ( .ip1(n2055), .ip2(n2054), .op(n2067) );
  inv_1 U2303 ( .ip(n2067), .op(n2060) );
  inv_1 U2304 ( .ip(n2056), .op(n2057) );
  nand2_1 U2305 ( .ip1(n2068), .ip2(n2059), .op(n2062) );
  nor2_1 U2306 ( .ip1(n2060), .ip2(n2062), .op(n2063) );
  nand2_1 U2307 ( .ip1(n2065), .ip2(n2066), .op(n2061) );
  nand2_1 U2308 ( .ip1(n2066), .ip2(n2065), .op(n2071) );
  nor3_1 U2309 ( .ip1(n2069), .ip2(n2068), .ip3(n2067), .op(n2070) );
  nand2_1 U2310 ( .ip1(n2071), .ip2(n2070), .op(n2072) );
  inv_1 U2311 ( .ip(n2074), .op(n2075) );
  nand2_1 U2312 ( .ip1(n2076), .ip2(n2075), .op(n2080) );
  nand2_1 U2313 ( .ip1(n2078), .ip2(\mult/storeQ [3]), .op(n2079) );
  nand2_1 U2314 ( .ip1(n2080), .ip2(n2079), .op(n622) );
  nand2_1 U2315 ( .ip1(n2082), .ip2(n2081), .op(n2090) );
  nor2_1 U2316 ( .ip1(n2084), .ip2(n2083), .op(n2088) );
  nor2_1 U2317 ( .ip1(n2086), .ip2(n2085), .op(n2087) );
  nor2_1 U2318 ( .ip1(n2088), .ip2(n2087), .op(n2089) );
  and2_1 U2319 ( .ip1(n2090), .ip2(n2089), .op(n2091) );
  nand2_1 U2320 ( .ip1(n2092), .ip2(n2091), .op(n2095) );
  nand2_1 U2321 ( .ip1(n2093), .ip2(\mult/storeQ [13]), .op(n2094) );
  nand2_1 U2322 ( .ip1(n2095), .ip2(n2094), .op(n612) );
  nand2_1 U2323 ( .ip1(n2137), .ip2(\mult/productQ [17]), .op(n2106) );
  and2_1 U2324 ( .ip1(n2097), .ip2(n2096), .op(n2103) );
  inv_1 U2325 ( .ip(n2098), .op(n2099) );
  nor2_1 U2326 ( .ip1(n2099), .ip2(n2126), .op(n2100) );
  nor2_1 U2327 ( .ip1(n2101), .ip2(n2100), .op(n2102) );
  nand2_1 U2328 ( .ip1(n2104), .ip2(n2151), .op(n2105) );
  nand2_1 U2329 ( .ip1(n2106), .ip2(n2105), .op(n576) );
  nand2_1 U2330 ( .ip1(n2137), .ip2(\mult/productQ [19]), .op(n2122) );
  and2_1 U2331 ( .ip1(n2109), .ip2(n2108), .op(n2119) );
  nand2_1 U2332 ( .ip1(n2110), .ip2(n2113), .op(n2112) );
  nand2_1 U2333 ( .ip1(n2112), .ip2(n2111), .op(n2117) );
  inv_1 U2334 ( .ip(n2113), .op(n2114) );
  nor2_1 U2335 ( .ip1(n2146), .ip2(n746), .op(n2116) );
  nor2_1 U2336 ( .ip1(n2117), .ip2(n2116), .op(n2118) );
  nand2_1 U2337 ( .ip1(n2122), .ip2(n2121), .op(n574) );
  and2_1 U2338 ( .ip1(n2125), .ip2(n2124), .op(n2134) );
  nand2_1 U2339 ( .ip1(n2145), .ip2(n2128), .op(n2127) );
  nand2_1 U2340 ( .ip1(n2141), .ip2(n2128), .op(n2130) );
  nand2_1 U2341 ( .ip1(n2135), .ip2(n1856), .op(n2136) );
  nand2_1 U2342 ( .ip1(n2137), .ip2(\mult/productQ [21]), .op(n2154) );
  nand2_1 U2343 ( .ip1(n2141), .ip2(n2144), .op(n2143) );
  nand2_1 U2344 ( .ip1(n2143), .ip2(n2142), .op(n2149) );
  nand2_1 U2345 ( .ip1(n2145), .ip2(n2144), .op(n2147) );
  nor2_1 U2346 ( .ip1(n2147), .ip2(n2146), .op(n2148) );
  nor2_1 U2347 ( .ip1(n2149), .ip2(n2148), .op(n2150) );
  nand2_1 U2348 ( .ip1(n2154), .ip2(n2153), .op(n572) );
  inv_1 U2349 ( .ip(\mult/state [0]), .op(n2155) );
  nor2_1 U2350 ( .ip1(\mult/state [1]), .ip2(n2155), .op(n2157) );
  not_ab_or_c_or_d U2351 ( .ip1(n2157), .ip2(\mult/counterQ [5]), .ip3(reset), 
        .ip4(n2156), .op(n632) );
  nand2_1 U2352 ( .ip1(n716), .ip2(doA[8]), .op(n2186) );
  nand2_1 U2353 ( .ip1(n716), .ip2(doA[6]), .op(n2185) );
  nand2_1 U2354 ( .ip1(n716), .ip2(doA[5]), .op(n2184) );
  nand2_1 U2355 ( .ip1(n716), .ip2(doB[7]), .op(n2170) );
  nand2_1 U2356 ( .ip1(n716), .ip2(doA[2]), .op(n2180) );
  nand2_1 U2357 ( .ip1(n716), .ip2(doA[1]), .op(n2181) );
  nand2_1 U2358 ( .ip1(n716), .ip2(doA[3]), .op(n2183) );
  nand2_1 U2359 ( .ip1(n716), .ip2(doA[4]), .op(n2182) );
  nand2_1 U2360 ( .ip1(n716), .ip2(doB[8]), .op(n2177) );
  nand2_1 U2361 ( .ip1(n716), .ip2(doB[15]), .op(n2164) );
  nand2_1 U2362 ( .ip1(n716), .ip2(doB[14]), .op(n2166) );
  nand2_1 U2363 ( .ip1(n716), .ip2(doB[3]), .op(n2171) );
  nand2_1 U2364 ( .ip1(n716), .ip2(doB[2]), .op(n2173) );
  nand2_1 U2365 ( .ip1(n716), .ip2(doB[1]), .op(n2174) );
  nand2_1 U2366 ( .ip1(n716), .ip2(doB[11]), .op(n2175) );
  nand2_1 U2367 ( .ip1(n716), .ip2(doB[13]), .op(n2165) );
  nand2_1 U2368 ( .ip1(n716), .ip2(doB[9]), .op(n2178) );
  nand2_1 U2369 ( .ip1(n716), .ip2(doB[10]), .op(n2176) );
  nand2_1 U2370 ( .ip1(n716), .ip2(doB[0]), .op(n2172) );
  nand2_1 U2371 ( .ip1(n716), .ip2(doB[5]), .op(n2169) );
  nand2_1 U2372 ( .ip1(n716), .ip2(doB[4]), .op(n2167) );
  nand2_1 U2373 ( .ip1(n716), .ip2(doB[6]), .op(n2168) );
  nand2_1 U2374 ( .ip1(n716), .ip2(doB[12]), .op(n2163) );
  nand2_1 U2375 ( .ip1(n716), .ip2(doA[0]), .op(n2179) );
  nand2_1 U2376 ( .ip1(n716), .ip2(doA[14]), .op(n2193) );
  nand2_1 U2377 ( .ip1(n716), .ip2(doA[9]), .op(n2188) );
  nand2_1 U2378 ( .ip1(n716), .ip2(doA[10]), .op(n2189) );
  nand2_1 U2379 ( .ip1(n716), .ip2(doA[7]), .op(n2187) );
  nand2_1 U2380 ( .ip1(n716), .ip2(doA[11]), .op(n2190) );
  nand2_1 U2381 ( .ip1(n716), .ip2(doA[12]), .op(n2191) );
  nand2_1 U2382 ( .ip1(n716), .ip2(doA[15]), .op(n2194) );
  nand2_1 U2383 ( .ip1(n716), .ip2(doA[13]), .op(n2192) );
  nand2_1 U2384 ( .ip1(n2228), .ip2(aBQ[0]), .op(n2201) );
  nand2_1 U2385 ( .ip1(n2225), .ip2(aAQ[0]), .op(n2217) );
  nand3_1 U2386 ( .ip1(n2228), .ip2(n2208), .ip3(aBQ[2]), .op(n2209) );
  nand3_1 U2387 ( .ip1(n2225), .ip2(n2224), .ip3(aAQ[2]), .op(n2226) );
  and2_1 U2388 ( .ip1(n2161), .ip2(aAQ[8]), .op(n16) );
  and2_1 U2389 ( .ip1(n2161), .ip2(aBQ[8]), .op(n17) );
  and2_1 U2390 ( .ip1(n2161), .ip2(aAQ[7]), .op(n15) );
  and2_1 U2391 ( .ip1(n2161), .ip2(aAQ[6]), .op(n14) );
  and2_1 U2392 ( .ip1(\nextState[0] ), .ip2(n2162), .op(n684) );
  mux2_1 U2393 ( .ip1(n2201), .ip2(n2205), .s(aBQ[1]), .op(n2202) );
  mux2_1 U2394 ( .ip1(n2206), .ip2(n2207), .s(aBQ[2]), .op(n2) );
  mux2_1 U2395 ( .ip1(n2225), .ip2(n2161), .s(aAQ[0]), .op(n8) );
  mux2_1 U2396 ( .ip1(n2217), .ip2(n2221), .s(aAQ[1]), .op(n2218) );
  mux2_1 U2397 ( .ip1(n2222), .ip2(n2223), .s(aAQ[2]), .op(n10) );
  mux2_1 U2398 ( .ip1(n2228), .ip2(n2161), .s(aBQ[0]), .op(n18) );
endmodule

