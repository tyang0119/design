`timescale 1ns / 1ps

module nopipe_tb();

    reg  [15:0] a;
    reg  [15:0] b;
    reg  clk;
    reg  reset;

    wire [15:0] product;

	//A = [ 1.25, 2.5, 2.5, 2, 3, 2, 1.25, 3.5, 4.5, 2]
	//B = [ 1.5, 1.5, 5, 2, 5, 3, 3.5, 5, 4, 3]


    mult DUT(
        .clk(clk),
        .reset(reset),
        .A(a),
        .B(b),
        .result(product)
        );

    initial
    begin
        $dumpfile("nopipe.vcd");
        $dumpvars(0, nopipe_tb);

        reset = 1;
        clk = 0;
        a = 0;
        b = 0;

        // 1
        #16
        reset = 0;
        a = 16'b0000000101000000;
        b = 16'b0000000110000000;
		// 2
        #1000
        a = 16'b0000001010000000;
        b = 16'b0000000110000000;

        // 3
        #1000		
        a = 16'b0000001010000000;
        b = 16'b0000010100000000;

        // 4
        #1000
        a = 16'b0000001000000000;
        b = 16'b0000001000000000;


        // 5
        #1000
        a = 16'b0000001100000000;
        b = 16'b0000010100000000;
		
        // 6
        #16
        a = 16'b0000001000000000;
        b = 16'b0000001100000000;


        // 7
        #1000
        a = 16'b0000000101000000;
        b = 16'b0000001110000000;

        // 8
        #1000
        a = 16'b0000001110000000;
        b = 16'b0000010100000000;

        // 9
        #1000
        a = 16'b0000010010000000;
        b = 16'b0000010000000000;


        // 10
        #1000
        a = 16'b0000001000000000;
        b = 16'b0000001100000000;
		
        $finish;
    end

    always 
        #10 clk = !clk;

endmodule