
module nopipe ( clk, reset, A, B, result, wrAddr );
  input [15:0] A;
  input [15:0] B;
  output [15:0] result;
  input [3:0] wrAddr;
  input clk, reset;
  wire   weB, N232, N233, N234, N235, N267, N268, N269, N270, N283, N284, N285,
         N286, N287, N288, N289, N290, N291, N292, N293, N294, N295, N296,
         N297, N298, N317, N318, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n530, n532, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n571, n572, n573, n574, n575, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n588, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957;
  wire   [8:0] aAQ;
  wire   [15:0] doA;
  wire   [8:0] aBQ;
  wire   [15:0] doB;
  wire   [15:0] result2;
  wire   [15:0] partialQ;
  wire   [1:0] state;
  wire   [15:0] counter2Q;
  wire   [15:0] counterQ;
  wire   [15:0] counterD;
  wire   [3:0] \mult/state ;
  wire   [6:0] \mult/counterQ ;
  wire   [31:0] \mult/productQ ;
  wire   [31:0] \mult/storeQ ;

  ramA rA ( .clk(clk), .we(weB), .a(aAQ), .di(A), .do(doA) );
  ramB rB ( .clk(clk), .we(weB), .a(aBQ), .di(B), .do(doB) );
  dp_1 \state_reg[1]  ( .ip(N318), .ck(clk), .q(state[1]) );
  dp_1 \partialQ_reg[8]  ( .ip(n449), .ck(clk), .q(partialQ[8]) );
  dp_1 \partialQ_reg[7]  ( .ip(n450), .ck(clk), .q(partialQ[7]) );
  dp_1 \partialQ_reg[6]  ( .ip(n451), .ck(clk), .q(partialQ[6]) );
  dp_1 \partialQ_reg[4]  ( .ip(n453), .ck(clk), .q(partialQ[4]) );
  dp_1 \partialQ_reg[3]  ( .ip(n454), .ck(clk), .q(partialQ[3]) );
  dp_1 \partialQ_reg[0]  ( .ip(n457), .ck(clk), .q(partialQ[0]) );
  dp_1 \counterQ_reg[0]  ( .ip(N267), .ck(clk), .q(counterQ[0]) );
  dp_1 \mult/state_reg[1]  ( .ip(n530), .ck(clk), .q(\mult/state [1]) );
  dp_1 \mult/state_reg[0]  ( .ip(n528), .ck(clk), .q(\mult/state [0]) );
  dp_1 \mult/counterQ_reg[5]  ( .ip(n527), .ck(clk), .q(\mult/counterQ [5]) );
  dp_1 \mult/storeQ_reg[17]  ( .ip(n504), .ck(clk), .q(\mult/storeQ [17]) );
  dp_1 \mult/storeQ_reg[21]  ( .ip(n500), .ck(clk), .q(\mult/storeQ [21]) );
  dp_1 \mult/storeQ_reg[13]  ( .ip(n508), .ck(clk), .q(\mult/storeQ [13]) );
  dp_1 \mult/storeQ_reg[7]  ( .ip(n514), .ck(clk), .q(\mult/storeQ [7]) );
  dp_1 \mult/storeQ_reg[23]  ( .ip(n498), .ck(clk), .q(\mult/storeQ [23]) );
  dp_1 \mult/storeQ_reg[15]  ( .ip(n506), .ck(clk), .q(\mult/storeQ [15]) );
  dp_1 \mult/storeQ_reg[6]  ( .ip(n515), .ck(clk), .q(\mult/storeQ [6]) );
  dp_1 \mult/storeQ_reg[22]  ( .ip(n499), .ck(clk), .q(\mult/storeQ [22]) );
  dp_1 \mult/storeQ_reg[14]  ( .ip(n507), .ck(clk), .q(\mult/storeQ [14]) );
  dp_1 \mult/storeQ_reg[2]  ( .ip(n519), .ck(clk), .q(\mult/storeQ [2]) );
  dp_1 \mult/storeQ_reg[18]  ( .ip(n503), .ck(clk), .q(\mult/storeQ [18]) );
  dp_1 \mult/storeQ_reg[10]  ( .ip(n511), .ck(clk), .q(\mult/storeQ [10]) );
  dp_1 \mult/storeQ_reg[4]  ( .ip(n517), .ck(clk), .q(\mult/storeQ [4]) );
  dp_1 \mult/storeQ_reg[20]  ( .ip(n501), .ck(clk), .q(\mult/storeQ [20]) );
  dp_1 \mult/storeQ_reg[12]  ( .ip(n509), .ck(clk), .q(\mult/storeQ [12]) );
  dp_1 \mult/storeQ_reg[16]  ( .ip(n505), .ck(clk), .q(\mult/storeQ [16]) );
  dp_1 \mult/productQ_reg[2]  ( .ip(n487), .ck(clk), .q(\mult/productQ [2]) );
  dp_1 \mult/productQ_reg[4]  ( .ip(n485), .ck(clk), .q(\mult/productQ [4]) );
  dp_1 \mult/productQ_reg[6]  ( .ip(n483), .ck(clk), .q(\mult/productQ [6]) );
  dp_1 \mult/productQ_reg[7]  ( .ip(n482), .ck(clk), .q(\mult/productQ [7]) );
  dp_1 \mult/productQ_reg[12]  ( .ip(n477), .ck(clk), .q(\mult/productQ [12])
         );
  dp_1 \mult/productQ_reg[13]  ( .ip(n476), .ck(clk), .q(\mult/productQ [13])
         );
  dp_1 \mult/productQ_reg[14]  ( .ip(n475), .ck(clk), .q(\mult/productQ [14])
         );
  dp_1 \mult/productQ_reg[15]  ( .ip(n474), .ck(clk), .q(\mult/productQ [15])
         );
  dp_1 \mult/productQ_reg[17]  ( .ip(n472), .ck(clk), .q(\mult/productQ [17])
         );
  dp_1 \mult/productQ_reg[20]  ( .ip(n469), .ck(clk), .q(\mult/productQ [20])
         );
  dp_1 \mult/productQ_reg[21]  ( .ip(n468), .ck(clk), .q(\mult/productQ [21])
         );
  dp_1 \mult/productQ_reg[22]  ( .ip(n467), .ck(clk), .q(\mult/productQ [22])
         );
  dp_1 \mult/productQ_reg[23]  ( .ip(n466), .ck(clk), .q(\mult/productQ [23])
         );
  lp_2 \mult/PRODUCT_reg[4]  ( .ck(n1173), .ip(\mult/productQ [12]), .q(
        result2[4]) );
  lp_2 \mult/PRODUCT_reg[5]  ( .ck(n1173), .ip(\mult/productQ [13]), .q(
        result2[5]) );
  lp_2 \mult/PRODUCT_reg[6]  ( .ck(n1173), .ip(\mult/productQ [14]), .q(
        result2[6]) );
  lp_2 \mult/PRODUCT_reg[8]  ( .ck(n1173), .ip(\mult/productQ [16]), .q(
        result2[8]) );
  lp_2 \mult/PRODUCT_reg[10]  ( .ck(n1173), .ip(\mult/productQ [18]), .q(
        result2[10]) );
  lp_2 \mult/PRODUCT_reg[11]  ( .ck(n1173), .ip(\mult/productQ [19]), .q(
        result2[11]) );
  lp_2 \mult/PRODUCT_reg[13]  ( .ck(n1173), .ip(\mult/productQ [21]), .q(
        result2[13]) );
  lp_2 \mult/PRODUCT_reg[14]  ( .ck(n1173), .ip(\mult/productQ [22]), .q(
        result2[14]) );
  dp_1 \aAQ_reg[0]  ( .ip(n18), .ck(clk), .q(aAQ[0]) );
  dp_1 \aBQ_reg[8]  ( .ip(n17), .ck(clk), .q(aBQ[8]) );
  dp_1 \aAQ_reg[8]  ( .ip(n16), .ck(clk), .q(aAQ[8]) );
  dp_1 \aAQ_reg[7]  ( .ip(n15), .ck(clk), .q(aAQ[7]) );
  dp_1 \aAQ_reg[6]  ( .ip(n14), .ck(clk), .q(aAQ[6]) );
  dp_1 \aAQ_reg[5]  ( .ip(n13), .ck(clk), .q(aAQ[5]) );
  dp_1 \aAQ_reg[3]  ( .ip(n11), .ck(clk), .q(aAQ[3]) );
  dp_1 \aAQ_reg[2]  ( .ip(n10), .ck(clk), .q(aAQ[2]) );
  dp_1 \aAQ_reg[1]  ( .ip(n9), .ck(clk), .q(aAQ[1]) );
  dp_1 \aBQ_reg[0]  ( .ip(n8), .ck(clk), .q(aBQ[0]) );
  dp_1 \aBQ_reg[1]  ( .ip(n7), .ck(clk), .q(aBQ[1]) );
  dp_1 \aBQ_reg[2]  ( .ip(n6), .ck(clk), .q(aBQ[2]) );
  dp_1 \aBQ_reg[3]  ( .ip(n5), .ck(clk), .q(aBQ[3]) );
  dp_1 \aBQ_reg[5]  ( .ip(n3), .ck(clk), .q(aBQ[5]) );
  dp_1 \aBQ_reg[6]  ( .ip(n2), .ck(clk), .q(aBQ[6]) );
  dp_1 \aBQ_reg[7]  ( .ip(n1), .ck(clk), .q(aBQ[7]) );
  inv_1 U607 ( .ip(n441), .op(weB) );
  dp_4 \mult/counterQ_reg[2]  ( .ip(n524), .ck(clk), .q(\mult/counterQ [2]) );
  lp_1 \mult/PRODUCT_reg[9]  ( .ck(n1173), .ip(\mult/productQ [17]), .q(
        result2[9]) );
  lp_1 \mult/PRODUCT_reg[1]  ( .ck(n1173), .ip(\mult/productQ [9]), .q(
        result2[1]) );
  dp_2 \mult/productQ_reg[18]  ( .ip(n471), .ck(clk), .q(\mult/productQ [18])
         );
  dp_2 \mult/storeQ_reg[5]  ( .ip(n516), .ck(clk), .q(\mult/storeQ [5]) );
  dp_2 \mult/productQ_reg[16]  ( .ip(n473), .ck(clk), .q(\mult/productQ [16])
         );
  dp_2 \mult/productQ_reg[1]  ( .ip(n488), .ck(clk), .q(\mult/productQ [1]) );
  dp_2 \mult/storeQ_reg[1]  ( .ip(n520), .ck(clk), .q(\mult/storeQ [1]) );
  dp_2 \mult/productQ_reg[10]  ( .ip(n479), .ck(clk), .q(\mult/productQ [10])
         );
  dp_2 \mult/productQ_reg[11]  ( .ip(n478), .ck(clk), .q(\mult/productQ [11])
         );
  dp_2 \mult/storeQ_reg[11]  ( .ip(n510), .ck(clk), .q(\mult/storeQ [11]) );
  dp_2 \mult/productQ_reg[0]  ( .ip(n489), .ck(clk), .q(\mult/productQ [0]) );
  dp_2 \mult/storeQ_reg[0]  ( .ip(n521), .ck(clk), .q(\mult/storeQ [0]) );
  dp_2 \mult/storeQ_reg[3]  ( .ip(n518), .ck(clk), .q(\mult/storeQ [3]) );
  dp_2 \mult/productQ_reg[3]  ( .ip(n486), .ck(clk), .q(\mult/productQ [3]) );
  dp_2 \mult/productQ_reg[19]  ( .ip(n470), .ck(clk), .q(\mult/productQ [19])
         );
  dp_2 \mult/storeQ_reg[19]  ( .ip(n502), .ck(clk), .q(\mult/storeQ [19]) );
  dp_2 \counterQ_reg[3]  ( .ip(N270), .ck(clk), .q(counterQ[3]) );
  dp_2 \mult/productQ_reg[8]  ( .ip(n481), .ck(clk), .q(\mult/productQ [8]) );
  dp_2 \mult/storeQ_reg[8]  ( .ip(n513), .ck(clk), .q(\mult/storeQ [8]) );
  dp_2 \counter2Q_reg[6]  ( .ip(N289), .ck(clk), .q(counter2Q[6]) );
  dp_2 \counter2Q_reg[2]  ( .ip(N285), .ck(clk), .q(counter2Q[2]) );
  dp_2 \counter2Q_reg[1]  ( .ip(N284), .ck(clk), .q(counter2Q[1]) );
  dp_2 \counter2Q_reg[5]  ( .ip(N288), .ck(clk), .q(counter2Q[5]) );
  dp_2 \counter2Q_reg[4]  ( .ip(N287), .ck(clk), .q(counter2Q[4]) );
  dp_2 \counter2Q_reg[9]  ( .ip(N292), .ck(clk), .q(counter2Q[9]) );
  dp_2 \counter2Q_reg[7]  ( .ip(N290), .ck(clk), .q(counter2Q[7]) );
  dp_1 \counterQ_reg[1]  ( .ip(N268), .ck(clk), .q(counterQ[1]) );
  dp_2 \mult/counterQ_reg[0]  ( .ip(n522), .ck(clk), .q(\mult/counterQ [0]) );
  dp_2 \partialQ_reg[15]  ( .ip(n442), .ck(clk), .q(partialQ[15]) );
  dp_2 \partialQ_reg[14]  ( .ip(n443), .ck(clk), .q(partialQ[14]) );
  dp_2 \mult/counterQ_reg[1]  ( .ip(n523), .ck(clk), .q(\mult/counterQ [1]) );
  dp_2 \state_reg[0]  ( .ip(N317), .ck(clk), .q(state[0]) );
  lp_1 \result_reg[14]  ( .ck(n532), .ip(partialQ[14]), .q(result[14]) );
  lp_1 \result_reg[11]  ( .ck(n532), .ip(partialQ[11]), .q(result[11]) );
  lp_1 \result_reg[0]  ( .ck(n532), .ip(partialQ[0]), .q(result[0]) );
  lp_1 \result_reg[15]  ( .ck(n532), .ip(partialQ[15]), .q(result[15]) );
  lp_1 \result_reg[6]  ( .ck(n532), .ip(partialQ[6]), .q(result[6]) );
  lp_1 \result_reg[12]  ( .ck(n532), .ip(partialQ[12]), .q(result[12]) );
  lp_1 \result_reg[8]  ( .ck(n532), .ip(partialQ[8]), .q(result[8]) );
  lp_1 \result_reg[7]  ( .ck(n532), .ip(partialQ[7]), .q(result[7]) );
  lp_1 \result_reg[4]  ( .ck(n532), .ip(partialQ[4]), .q(result[4]) );
  lp_1 \result_reg[2]  ( .ck(n532), .ip(partialQ[2]), .q(result[2]) );
  lp_1 \result_reg[5]  ( .ck(n532), .ip(partialQ[5]), .q(result[5]) );
  lp_1 \result_reg[13]  ( .ck(n532), .ip(partialQ[13]), .q(result[13]) );
  lp_1 \result_reg[10]  ( .ck(n532), .ip(partialQ[10]), .q(result[10]) );
  lp_1 \result_reg[9]  ( .ck(n532), .ip(partialQ[9]), .q(result[9]) );
  lp_1 \result_reg[3]  ( .ck(n532), .ip(partialQ[3]), .q(result[3]) );
  lp_1 \result_reg[1]  ( .ck(n532), .ip(partialQ[1]), .q(result[1]) );
  lp_1 \mult/PRODUCT_reg[3]  ( .ck(n1173), .ip(\mult/productQ [11]), .q(
        result2[3]) );
  lp_1 \mult/PRODUCT_reg[0]  ( .ck(n1173), .ip(\mult/productQ [8]), .q(
        result2[0]) );
  dp_2 \mult/productQ_reg[5]  ( .ip(n484), .ck(clk), .q(\mult/productQ [5]) );
  dp_2 \counter2Q_reg[14]  ( .ip(N297), .ck(clk), .q(counter2Q[14]) );
  dp_2 \mult/storeQ_reg[9]  ( .ip(n512), .ck(clk), .q(\mult/storeQ [9]) );
  dp_2 \mult/productQ_reg[9]  ( .ip(n480), .ck(clk), .q(\mult/productQ [9]) );
  dp_2 \counter2Q_reg[8]  ( .ip(N291), .ck(clk), .q(counter2Q[8]) );
  dp_2 \counter2Q_reg[0]  ( .ip(N283), .ck(clk), .q(counter2Q[0]) );
  dp_2 \counter2Q_reg[15]  ( .ip(N298), .ck(clk), .q(counter2Q[15]) );
  dp_2 \counter2Q_reg[13]  ( .ip(N296), .ck(clk), .q(counter2Q[13]) );
  dp_2 \counter2Q_reg[11]  ( .ip(N294), .ck(clk), .q(counter2Q[11]) );
  dp_2 \counter2Q_reg[12]  ( .ip(N295), .ck(clk), .q(counter2Q[12]) );
  dp_2 \partialQ_reg[12]  ( .ip(n445), .ck(clk), .q(partialQ[12]) );
  dksp_1 \mult/counterQ_reg[4]  ( .ip(n526), .sb(1'b1), .ck(clk), .q(n671), 
        .qb() );
  dp_2 \partialQ_reg[1]  ( .ip(n456), .ck(clk), .q(partialQ[1]) );
  dp_2 \partialQ_reg[5]  ( .ip(n452), .ck(clk), .q(partialQ[5]) );
  dp_2 \partialQ_reg[13]  ( .ip(n444), .ck(clk), .q(partialQ[13]) );
  dp_2 \partialQ_reg[2]  ( .ip(n455), .ck(clk), .q(partialQ[2]) );
  lp_1 \mult/PRODUCT_reg[12]  ( .ck(n1849), .ip(\mult/productQ [20]), .q(
        result2[12]) );
  dp_2 \partialQ_reg[9]  ( .ip(n448), .ck(clk), .q(partialQ[9]) );
  dp_4 \mult/counterQ_reg[3]  ( .ip(n525), .ck(clk), .q(\mult/counterQ [3]) );
  lp_1 \counterD_reg[0]  ( .ck(n1957), .ip(N232), .q(counterD[0]) );
  lp_1 \counterD_reg[1]  ( .ck(n1957), .ip(N233), .q(counterD[1]) );
  lp_1 \counterD_reg[2]  ( .ck(n1957), .ip(N234), .q(counterD[2]) );
  lp_1 \counterD_reg[3]  ( .ck(n1957), .ip(N235), .q(counterD[3]) );
  dp_1 \counter2Q_reg[10]  ( .ip(N293), .ck(clk), .q(counter2Q[10]) );
  dp_2 \counterQ_reg[2]  ( .ip(N269), .ck(clk), .q(counterQ[2]) );
  dp_1 \counter2Q_reg[3]  ( .ip(N286), .ck(clk), .q(counter2Q[3]) );
  dp_2 \partialQ_reg[11]  ( .ip(n446), .ck(clk), .q(partialQ[11]) );
  lp_1 \mult/PRODUCT_reg[7]  ( .ck(n1173), .ip(\mult/productQ [15]), .q(
        result2[7]) );
  dp_2 \partialQ_reg[10]  ( .ip(n447), .ck(clk), .q(partialQ[10]) );
  lp_1 \mult/PRODUCT_reg[2]  ( .ck(n1173), .ip(\mult/productQ [10]), .q(
        result2[2]) );
  lp_1 \mult/PRODUCT_reg[15]  ( .ck(n1173), .ip(\mult/productQ [23]), .q(
        result2[15]) );
  dp_1 \aAQ_reg[4]  ( .ip(n12), .ck(clk), .q(aAQ[4]) );
  dp_1 \aBQ_reg[4]  ( .ip(n4), .ck(clk), .q(aBQ[4]) );
  inv_2 U608 ( .ip(n710), .op(n1833) );
  inv_1 U609 ( .ip(aBQ[3]), .op(n1900) );
  buf_2 U610 ( .ip(n999), .op(n1767) );
  buf_4 U611 ( .ip(n955), .op(n1470) );
  nor2_2 U612 ( .ip1(n1821), .ip2(n1164), .op(n1165) );
  nor2_1 U613 ( .ip1(n946), .ip2(n1845), .op(n947) );
  nor2_2 U614 ( .ip1(n1574), .ip2(n1008), .op(n1803) );
  mux2_2 U615 ( .ip1(n1923), .ip2(n1922), .s(aBQ[1]), .op(n7) );
  nand2_1 U616 ( .ip1(n1811), .ip2(n1783), .op(n1813) );
  buf_4 U617 ( .ip(n1022), .op(n1480) );
  buf_4 U618 ( .ip(n1022), .op(n1519) );
  nand2_1 U619 ( .ip1(n1579), .ip2(n1783), .op(n1581) );
  nor2_2 U620 ( .ip1(n995), .ip2(n994), .op(n1002) );
  mux2_2 U621 ( .ip1(n1906), .ip2(n1905), .s(aBQ[6]), .op(n2) );
  nor2_1 U622 ( .ip1(n1927), .ip2(n1845), .op(n1838) );
  nand4_1 U623 ( .ip1(n1848), .ip2(\mult/counterQ [2]), .ip3(n1175), .ip4(
        doB[4]), .op(n1846) );
  inv_1 U624 ( .ip(n1851), .op(n1848) );
  nand2_1 U625 ( .ip1(n1274), .ip2(n1833), .op(n1276) );
  nand2_4 U626 ( .ip1(n1002), .ip2(n1001), .op(n1802) );
  nand3_2 U627 ( .ip1(n902), .ip2(n901), .ip3(n900), .op(n1036) );
  nor2_4 U628 ( .ip1(n1349), .ip2(n1892), .op(n1469) );
  nand2_1 U629 ( .ip1(n736), .ip2(n735), .op(n645) );
  inv_2 U630 ( .ip(n1620), .op(n1145) );
  nand2_2 U631 ( .ip1(n1825), .ip2(partialQ[15]), .op(n1644) );
  nand2_1 U632 ( .ip1(n794), .ip2(n599), .op(n796) );
  or2_2 U633 ( .ip1(n777), .ip2(n778), .op(n794) );
  nand2_2 U634 ( .ip1(n626), .ip2(n882), .op(n880) );
  nand2_2 U635 ( .ip1(n624), .ip2(n610), .op(n626) );
  inv_1 U636 ( .ip(result2[5]), .op(n719) );
  inv_1 U637 ( .ip(n898), .op(n901) );
  nor2_1 U638 ( .ip1(n1264), .ip2(n765), .op(n731) );
  nor2_1 U639 ( .ip1(n1040), .ip2(n1039), .op(n1041) );
  inv_1 U640 ( .ip(n671), .op(n1034) );
  inv_1 U641 ( .ip(n1635), .op(n1135) );
  nor2_1 U642 ( .ip1(n1317), .ip2(n1316), .op(n1386) );
  inv_1 U643 ( .ip(n1854), .op(n1847) );
  nand2_1 U644 ( .ip1(n1824), .ip2(n1833), .op(n1827) );
  or2_1 U645 ( .ip1(n539), .ip2(n1448), .op(n535) );
  or2_1 U646 ( .ip1(n539), .ip2(n1475), .op(n536) );
  or2_1 U647 ( .ip1(n539), .ip2(n1460), .op(n537) );
  xnor2_2 U648 ( .ip1(n1071), .ip2(n1068), .op(n538) );
  or2_1 U649 ( .ip1(\mult/counterQ [3]), .ip2(n671), .op(n539) );
  nand2_1 U650 ( .ip1(n540), .ip2(n1151), .op(n1157) );
  inv_1 U651 ( .ip(n1149), .op(n540) );
  nand2_1 U652 ( .ip1(n1130), .ip2(n619), .op(n1149) );
  nand2_1 U653 ( .ip1(n1615), .ip2(n619), .op(n1632) );
  nor2_1 U654 ( .ip1(n1264), .ip2(n764), .op(n544) );
  nor2_1 U655 ( .ip1(n543), .ip2(n541), .op(n1452) );
  nand2_1 U656 ( .ip1(n542), .ip2(n535), .op(n541) );
  nand2_1 U657 ( .ip1(n1451), .ip2(\mult/counterQ [3]), .op(n542) );
  nor2_1 U658 ( .ip1(n1449), .ip2(n1506), .op(n543) );
  nand2_1 U659 ( .ip1(n545), .ip2(n544), .op(n639) );
  inv_1 U660 ( .ip(n638), .op(n545) );
  nand2_1 U661 ( .ip1(n1486), .ip2(n546), .op(n795) );
  nand2_1 U662 ( .ip1(n840), .ip2(n718), .op(n546) );
  inv_1 U663 ( .ip(n547), .op(n661) );
  nand3_1 U664 ( .ip1(n1633), .ip2(n1833), .ip3(n1634), .op(n547) );
  or2_1 U665 ( .ip1(n1626), .ip2(partialQ[15]), .op(n1634) );
  and2_1 U666 ( .ip1(result2[9]), .ip2(n733), .op(n803) );
  or2_1 U667 ( .ip1(n800), .ip2(n1624), .op(n582) );
  nand2_1 U668 ( .ip1(n1401), .ip2(n655), .op(n1356) );
  nand2_1 U669 ( .ip1(n1814), .ip2(n727), .op(n742) );
  inv_1 U670 ( .ip(n549), .op(n649) );
  nand3_1 U671 ( .ip1(n1868), .ip2(n1869), .ip3(\mult/counterQ [3]), .op(n549)
         );
  and2_1 U672 ( .ip1(n733), .ip2(result2[4]), .op(n746) );
  nand2_1 U673 ( .ip1(n1614), .ip2(n1557), .op(n605) );
  nand2_1 U674 ( .ip1(n618), .ip2(n871), .op(n1614) );
  inv_1 U675 ( .ip(n550), .op(n652) );
  nand2_1 U676 ( .ip1(n1034), .ip2(n1036), .op(n550) );
  nand2_1 U677 ( .ip1(n1518), .ip2(n551), .op(n1482) );
  nor2_1 U678 ( .ip1(n552), .ip2(n1477), .op(n551) );
  nand2_1 U679 ( .ip1(n553), .ip2(n536), .op(n552) );
  nand2_1 U680 ( .ip1(n1478), .ip2(\mult/counterQ [3]), .op(n553) );
  nand3_1 U681 ( .ip1(n1571), .ip2(n554), .ip3(n555), .op(n445) );
  nand2_1 U682 ( .ip1(n1562), .ip2(n1561), .op(n554) );
  nand2_1 U683 ( .ip1(n1568), .ip2(n1565), .op(n555) );
  inv_1 U684 ( .ip(n848), .op(n1159) );
  nand2_1 U685 ( .ip1(n853), .ip2(n852), .op(n848) );
  nand2_1 U686 ( .ip1(n608), .ip2(n556), .op(n1610) );
  inv_1 U687 ( .ip(n557), .op(n556) );
  nand2_1 U688 ( .ip1(n1595), .ip2(n1589), .op(n557) );
  nand2_1 U689 ( .ip1(n559), .ip2(n558), .op(n638) );
  inv_1 U690 ( .ip(n765), .op(n558) );
  inv_1 U691 ( .ip(n800), .op(n559) );
  nand2_1 U692 ( .ip1(n1518), .ip2(n560), .op(n1466) );
  nor2_1 U693 ( .ip1(n561), .ip2(n1462), .op(n560) );
  nand2_1 U694 ( .ip1(n562), .ip2(n537), .op(n561) );
  nand2_1 U695 ( .ip1(n1463), .ip2(\mult/counterQ [3]), .op(n562) );
  nand2_1 U696 ( .ip1(n563), .ip2(n1520), .op(n500) );
  nand2_1 U697 ( .ip1(n564), .ip2(n1518), .op(n563) );
  inv_1 U698 ( .ip(n565), .op(n564) );
  nand2_1 U699 ( .ip1(n1517), .ip2(n1516), .op(n565) );
  nand2_1 U700 ( .ip1(n709), .ip2(n711), .op(n712) );
  and2_1 U701 ( .ip1(n782), .ip2(n781), .op(n566) );
  nand2_2 U702 ( .ip1(n830), .ip2(n1544), .op(n1905) );
  nand2_2 U703 ( .ip1(n824), .ip2(n1544), .op(n1922) );
  nor2_1 U704 ( .ip1(n789), .ip2(n639), .op(n1295) );
  inv_1 U705 ( .ip(n1443), .op(n1511) );
  nand2_1 U706 ( .ip1(n1619), .ip2(n1612), .op(n1616) );
  nand2_2 U707 ( .ip1(n1525), .ip2(n749), .op(n750) );
  nand2_1 U708 ( .ip1(n739), .ip2(n726), .op(n730) );
  inv_2 U709 ( .ip(n591), .op(n863) );
  nor2_4 U710 ( .ip1(n851), .ip2(n850), .op(n852) );
  xnor2_1 U711 ( .ip1(n600), .ip2(n1809), .op(n1811) );
  xnor2_1 U712 ( .ip1(n602), .ip2(n1578), .op(n1579) );
  inv_2 U713 ( .ip(n569), .op(n567) );
  inv_2 U714 ( .ip(n761), .op(n768) );
  nor2_2 U715 ( .ip1(aAQ[1]), .ip2(n1945), .op(n1845) );
  nand2_1 U716 ( .ip1(n727), .ip2(n1814), .op(n729) );
  nor2_1 U717 ( .ip1(n665), .ip2(n1261), .op(n732) );
  inv_2 U718 ( .ip(n640), .op(n568) );
  inv_1 U719 ( .ip(result2[1]), .op(n734) );
  nand2_1 U720 ( .ip1(result2[12]), .ip2(n1622), .op(n861) );
  and2_1 U721 ( .ip1(n988), .ip2(n1705), .op(n989) );
  nor2_1 U722 ( .ip1(n1009), .ip2(n1803), .op(n1010) );
  nand2_1 U723 ( .ip1(n931), .ip2(n930), .op(n1371) );
  inv_2 U724 ( .ip(n710), .op(n711) );
  nand2_1 U725 ( .ip1(n992), .ip2(n991), .op(n1499) );
  inv_1 U726 ( .ip(n1225), .op(n571) );
  nor2_1 U727 ( .ip1(n1900), .ip2(n1860), .op(n1861) );
  inv_1 U728 ( .ip(\mult/productQ [1]), .op(n915) );
  inv_2 U729 ( .ip(aAQ[3]), .op(n1859) );
  nor3_2 U730 ( .ip1(aBQ[2]), .ip2(aBQ[1]), .ip3(aBQ[0]), .op(n1860) );
  inv_1 U731 ( .ip(\mult/storeQ [1]), .op(n914) );
  nor3_4 U732 ( .ip1(aBQ[4]), .ip2(aBQ[6]), .ip3(aBQ[5]), .op(n1898) );
  and2_1 U733 ( .ip1(state[0]), .ip2(n1181), .op(n684) );
  inv_1 U734 ( .ip(partialQ[9]), .op(n806) );
  nor2_1 U735 ( .ip1(aBQ[8]), .ip2(aAQ[5]), .op(n1857) );
  nor2_1 U736 ( .ip1(aAQ[7]), .ip2(aAQ[8]), .op(n1856) );
  nand2_1 U737 ( .ip1(n1168), .ip2(n1167), .op(n455) );
  nor2_1 U738 ( .ip1(n1628), .ip2(n1627), .op(n1629) );
  nand2_1 U739 ( .ip1(n943), .ip2(n942), .op(n480) );
  nand2_1 U740 ( .ip1(n845), .ip2(n567), .op(n653) );
  inv_1 U741 ( .ip(n865), .op(n881) );
  inv_1 U742 ( .ip(n1616), .op(n1617) );
  nand2_1 U743 ( .ip1(n1295), .ip2(n768), .op(n771) );
  inv_1 U744 ( .ip(n1263), .op(n1787) );
  nor2_1 U745 ( .ip1(n748), .ip2(n596), .op(n749) );
  nor2_1 U746 ( .ip1(n1529), .ip2(n1528), .op(n1532) );
  inv_2 U747 ( .ip(n1619), .op(n1134) );
  inv_1 U748 ( .ip(n634), .op(n1591) );
  inv_2 U749 ( .ip(n1549), .op(n569) );
  nand2_2 U750 ( .ip1(n730), .ip2(n729), .op(n761) );
  inv_1 U751 ( .ip(n796), .op(n797) );
  nand2_1 U752 ( .ip1(n732), .ip2(n863), .op(n737) );
  inv_1 U753 ( .ip(n1788), .op(n736) );
  nand2_1 U754 ( .ip1(n1131), .ip2(n762), .op(n1788) );
  inv_1 U755 ( .ip(n1261), .op(n1262) );
  nor2_1 U756 ( .ip1(n790), .ip2(n789), .op(n791) );
  nand2_1 U757 ( .ip1(n623), .ip2(n1268), .op(n830) );
  nand2_1 U758 ( .ip1(n1000), .ip2(n999), .op(n1001) );
  nand2_2 U759 ( .ip1(n1135), .ip2(n636), .op(n642) );
  inv_2 U760 ( .ip(n582), .op(n1138) );
  inv_2 U761 ( .ip(n727), .op(n741) );
  inv_1 U762 ( .ip(n861), .op(n862) );
  nor2_1 U763 ( .ip1(n1028), .ip2(n1027), .op(n1423) );
  inv_1 U764 ( .ip(n934), .op(n935) );
  inv_1 U765 ( .ip(result2[8]), .op(n625) );
  nor2_1 U766 ( .ip1(n1200), .ip2(n1178), .op(n1255) );
  nand2_1 U767 ( .ip1(n927), .ip2(n933), .op(n934) );
  xor2_2 U768 ( .ip1(n1668), .ip2(n1667), .op(n648) );
  nand4_1 U769 ( .ip1(n1430), .ip2(n1429), .ip3(n1428), .ip4(n1427), .op(n1442) );
  xnor2_1 U770 ( .ip1(n1247), .ip2(counterQ[3]), .op(n1248) );
  nand2_1 U771 ( .ip1(n1330), .ip2(n1329), .op(n1461) );
  nand4_1 U772 ( .ip1(n1397), .ip2(n1396), .ip3(n1395), .ip4(n1394), .op(n1467) );
  and2_1 U773 ( .ip1(n1340), .ip2(n1339), .op(n1341) );
  xnor2_1 U774 ( .ip1(n1234), .ip2(n616), .op(n1235) );
  nand3_1 U775 ( .ip1(n1334), .ip2(n1333), .ip3(n1881), .op(n1449) );
  nand4_1 U776 ( .ip1(n1437), .ip2(n1436), .ip3(n1435), .ip4(n1434), .op(n1455) );
  xnor2_1 U777 ( .ip1(n1230), .ip2(n1233), .op(n1231) );
  inv_1 U778 ( .ip(n1184), .op(n1668) );
  nand2_1 U779 ( .ip1(n656), .ip2(n897), .op(n898) );
  xnor2_1 U780 ( .ip1(n1251), .ip2(n1245), .op(n1252) );
  nand2_1 U781 ( .ip1(n932), .ip2(n1371), .op(n933) );
  nand2_1 U782 ( .ip1(n1091), .ip2(n1090), .op(n1097) );
  and2_1 U783 ( .ip1(n926), .ip2(n1369), .op(n927) );
  nor2_1 U784 ( .ip1(n1182), .ip2(n1229), .op(n1184) );
  nand2_1 U785 ( .ip1(n1499), .ip2(n997), .op(n993) );
  nor2_1 U786 ( .ip1(n1216), .ip2(n1215), .op(n1680) );
  nor3_2 U787 ( .ip1(n441), .ip2(n688), .ip3(n1828), .op(n689) );
  mux2_1 U788 ( .ip1(n1885), .ip2(n1884), .s(n1853), .op(n1406) );
  nor3_2 U789 ( .ip1(aBQ[7]), .ip2(n1862), .ip3(n1861), .op(n1899) );
  nor2_1 U790 ( .ip1(n1110), .ip2(n1114), .op(n1078) );
  nor2_1 U791 ( .ip1(n671), .ip2(n1035), .op(n1037) );
  mux2_1 U792 ( .ip1(n1877), .ip2(n1876), .s(n1853), .op(n1342) );
  nor2_1 U793 ( .ip1(n1056), .ip2(n918), .op(n919) );
  buf_1 U794 ( .ip(n1849), .op(n1173) );
  mux2_1 U795 ( .ip1(n1879), .ip2(n1878), .s(n1853), .op(n1318) );
  mux2_1 U796 ( .ip1(n1875), .ip2(n1874), .s(n1853), .op(n1316) );
  mux2_1 U797 ( .ip1(doA[4]), .ip2(doA[3]), .s(n1853), .op(n1886) );
  nand2_1 U798 ( .ip1(n1693), .ip2(n929), .op(n930) );
  and2_1 U799 ( .ip1(n1244), .ip2(counterQ[0]), .op(n1245) );
  nand3_1 U800 ( .ip1(n1857), .ip2(n1856), .ip3(n1855), .op(n1828) );
  inv_1 U801 ( .ip(n1698), .op(n929) );
  inv_1 U802 ( .ip(n806), .op(n805) );
  inv_1 U803 ( .ip(n1789), .op(n735) );
  inv_1 U804 ( .ip(n1195), .op(n903) );
  nor2_1 U805 ( .ip1(n1096), .ip2(n1095), .op(n1100) );
  inv_1 U806 ( .ip(n1076), .op(n1114) );
  inv_1 U807 ( .ip(n615), .op(n616) );
  nor2_1 U808 ( .ip1(n1934), .ip2(n1933), .op(n1942) );
  inv_1 U809 ( .ip(n1512), .op(n1035) );
  nor2_1 U810 ( .ip1(n1361), .ip2(n1057), .op(n918) );
  nand2_1 U811 ( .ip1(n922), .ip2(n921), .op(n1374) );
  xnor2_1 U812 ( .ip1(counterQ[0]), .ip2(n1253), .op(n1254) );
  nand2_2 U813 ( .ip1(n684), .ip2(n1586), .op(n710) );
  nand2_1 U814 ( .ip1(n924), .ip2(n923), .op(n1370) );
  buf_1 U815 ( .ip(partialQ[5]), .op(n787) );
  inv_2 U816 ( .ip(counterQ[2]), .op(n681) );
  inv_1 U817 ( .ip(partialQ[0]), .op(n1264) );
  inv_1 U818 ( .ip(partialQ[1]), .op(n1789) );
  inv_1 U819 ( .ip(partialQ[2]), .op(n726) );
  buf_1 U820 ( .ip(partialQ[15]), .op(n1625) );
  inv_2 U821 ( .ip(partialQ[14]), .op(n1133) );
  inv_1 U822 ( .ip(partialQ[6]), .op(n1486) );
  nand2_1 U823 ( .ip1(\mult/productQ [4]), .ip2(\mult/storeQ [4]), .op(n1698)
         );
  inv_1 U824 ( .ip(partialQ[11]), .op(n1594) );
  or2_1 U825 ( .ip1(\mult/storeQ [5]), .ip2(\mult/productQ [5]), .op(n1693) );
  inv_1 U826 ( .ip(aAQ[2]), .op(n1930) );
  nand2_1 U827 ( .ip1(aAQ[2]), .ip2(aAQ[0]), .op(n1934) );
  nand2_1 U828 ( .ip1(aAQ[3]), .ip2(aAQ[1]), .op(n1933) );
  inv_1 U829 ( .ip(aAQ[7]), .op(n1950) );
  inv_1 U830 ( .ip(aBQ[7]), .op(n1954) );
  inv_2 U831 ( .ip(\mult/counterQ [3]), .op(n1512) );
  inv_1 U832 ( .ip(aBQ[2]), .op(n1917) );
  nor3_4 U833 ( .ip1(aAQ[0]), .ip2(aAQ[2]), .ip3(aAQ[1]), .op(n1858) );
  inv_2 U834 ( .ip(n802), .op(n789) );
  nand2_2 U835 ( .ip1(n572), .ip2(n705), .op(n706) );
  nor2_2 U836 ( .ip1(counter2Q[9]), .ip2(counter2Q[13]), .op(n572) );
  nor2_2 U837 ( .ip1(counter2Q[7]), .ip2(counter2Q[9]), .op(n673) );
  nand4_1 U838 ( .ip1(n853), .ip2(n852), .ip3(result2[10]), .ip4(n733), .op(
        n857) );
  nor2_2 U839 ( .ip1(counter2Q[11]), .ip2(counter2Q[13]), .op(n674) );
  nand2_2 U840 ( .ip1(n612), .ip2(n849), .op(n859) );
  nand2_2 U841 ( .ip1(counter2Q[1]), .ip2(counter2Q[2]), .op(n678) );
  nor2_2 U842 ( .ip1(counter2Q[4]), .ip2(counter2Q[8]), .op(n672) );
  buf_1 U843 ( .ip(n1774), .op(n573) );
  nor3_1 U844 ( .ip1(n611), .ip2(n569), .ip3(n868), .op(n869) );
  nand2_1 U845 ( .ip1(n1587), .ip2(n856), .op(n611) );
  nor2_2 U846 ( .ip1(n895), .ip2(n894), .op(n902) );
  nand2_1 U847 ( .ip1(n1732), .ip2(n574), .op(n476) );
  nand2_4 U848 ( .ip1(n1731), .ip2(n1810), .op(n574) );
  nand2_1 U849 ( .ip1(n1742), .ip2(n575), .op(n475) );
  nand2_4 U850 ( .ip1(n1741), .ip2(n1810), .op(n575) );
  nand2_2 U851 ( .ip1(n892), .ip2(n1873), .op(n907) );
  nand3_1 U852 ( .ip1(doB[1]), .ip2(n1870), .ip3(n1892), .op(n1872) );
  nor2_2 U853 ( .ip1(n1175), .ip2(\mult/counterQ [1]), .op(n1870) );
  nand2_1 U854 ( .ip1(n1585), .ip2(n577), .op(n471) );
  nand2_2 U855 ( .ip1(n1584), .ip2(n1810), .op(n577) );
  nand2_2 U856 ( .ip1(n853), .ip2(n852), .op(n620) );
  buf_1 U857 ( .ip(counter2Q[7]), .op(n578) );
  buf_1 U858 ( .ip(counter2Q[11]), .op(n579) );
  inv_1 U859 ( .ip(n580), .op(n1556) );
  nand2_1 U860 ( .ip1(n621), .ip2(n581), .op(n580) );
  nand2_1 U861 ( .ip1(n626), .ip2(n1550), .op(n581) );
  inv_4 U862 ( .ip(n1624), .op(n802) );
  nand2_4 U863 ( .ip1(n708), .ip2(n707), .op(n1624) );
  nand2_2 U864 ( .ip1(n1292), .ip2(n1549), .op(n583) );
  nand2_1 U865 ( .ip1(n1292), .ip2(n1549), .op(n846) );
  nor2_2 U866 ( .ip1(n586), .ip2(n1623), .op(n1626) );
  inv_1 U867 ( .ip(n1657), .op(n584) );
  inv_1 U868 ( .ip(n1223), .op(n585) );
  inv_1 U869 ( .ip(n802), .op(n586) );
  or2_2 U870 ( .ip1(n1283), .ip2(n1506), .op(n1518) );
  nand2_2 U871 ( .ip1(n967), .ip2(n966), .op(n974) );
  nand2_2 U872 ( .ip1(n725), .ip2(result2[7]), .op(n716) );
  inv_2 U873 ( .ip(n974), .op(n1042) );
  nand2_1 U874 ( .ip1(n840), .ip2(n718), .op(n598) );
  nand2_1 U875 ( .ip1(n683), .ip2(counterQ[3]), .op(n588) );
  nand2_1 U876 ( .ip1(n1159), .ip2(n590), .op(n744) );
  and2_1 U877 ( .ip1(n741), .ip2(partialQ[3]), .op(n590) );
  inv_1 U878 ( .ip(n802), .op(n591) );
  nand2_1 U879 ( .ip1(n1026), .ip2(n1025), .op(n592) );
  nor2_1 U880 ( .ip1(n592), .ip2(n593), .op(n651) );
  or2_1 U881 ( .ip1(n594), .ip2(n1028), .op(n593) );
  inv_1 U882 ( .ip(n1045), .op(n594) );
  inv_4 U883 ( .ip(\mult/counterQ [2]), .op(n1892) );
  nor2_4 U884 ( .ip1(\mult/counterQ [2]), .ip2(n1445), .op(n1850) );
  ab_or_c_or_d U885 ( .ip1(n1880), .ip2(doB[12]), .ip3(n1843), .ip4(n1839), 
        .op(n595) );
  mux2_2 U886 ( .ip1(n1200), .ip2(n966), .s(n1847), .op(n522) );
  nand2_2 U887 ( .ip1(n1899), .ip2(n689), .op(n690) );
  xnor2_2 U888 ( .ip1(n1818), .ip2(n1823), .op(n1824) );
  nand2_1 U889 ( .ip1(n1527), .ip2(n1272), .op(n596) );
  nand2_2 U890 ( .ip1(n1522), .ip2(n747), .op(n1272) );
  nand3_2 U891 ( .ip1(n1160), .ip2(n840), .ip3(n742), .op(n743) );
  nand2_1 U892 ( .ip1(n784), .ip2(n718), .op(n597) );
  nand2_1 U893 ( .ip1(n1159), .ip2(n718), .op(n773) );
  nand2_1 U894 ( .ip1(n1486), .ip2(n598), .op(n599) );
  or2_1 U895 ( .ip1(n1798), .ip2(n1797), .op(n600) );
  nand2_2 U896 ( .ip1(n583), .ip2(n845), .op(n613) );
  xnor2_1 U897 ( .ip1(n601), .ip2(n1583), .op(n1584) );
  or2_1 U898 ( .ip1(n1804), .ip2(n1806), .op(n601) );
  nand2_2 U899 ( .ip1(n1587), .ip2(n856), .op(n1128) );
  or2_1 U900 ( .ip1(n1575), .ip2(n1574), .op(n602) );
  inv_1 U901 ( .ip(n770), .op(n603) );
  buf_1 U902 ( .ip(n1535), .op(n604) );
  nand2_1 U903 ( .ip1(n608), .ip2(n1589), .op(n606) );
  inv_1 U904 ( .ip(n1508), .op(n607) );
  inv_1 U905 ( .ip(n1621), .op(n1638) );
  inv_1 U906 ( .ip(n1563), .op(n1564) );
  nand2_2 U907 ( .ip1(n784), .ip2(n783), .op(n785) );
  nand2_1 U908 ( .ip1(n872), .ip2(n871), .op(n608) );
  nand2_2 U909 ( .ip1(n776), .ip2(n1293), .op(n609) );
  nand2_1 U910 ( .ip1(n776), .ip2(n1293), .op(n610) );
  nand2_1 U911 ( .ip1(n776), .ip2(n1293), .op(n871) );
  inv_1 U912 ( .ip(n848), .op(n612) );
  nand2_4 U913 ( .ip1(\mult/counterQ [2]), .ip2(n893), .op(n1443) );
  nand2_4 U914 ( .ip1(n682), .ip2(n681), .op(n683) );
  inv_2 U915 ( .ip(counterQ[1]), .op(n682) );
  nand2_2 U916 ( .ip1(n1519), .ip2(\mult/storeQ [19]), .op(n1353) );
  nand2_2 U917 ( .ip1(n1036), .ip2(n595), .op(n949) );
  nand2_1 U918 ( .ip1(n845), .ip2(n846), .op(n614) );
  nand2_2 U919 ( .ip1(n805), .ip2(n804), .op(n845) );
  inv_1 U920 ( .ip(counter2Q[3]), .op(n615) );
  inv_1 U921 ( .ip(n1204), .op(n617) );
  and2_1 U922 ( .ip1(n722), .ip2(n1487), .op(n723) );
  inv_2 U923 ( .ip(n1291), .op(n618) );
  inv_1 U924 ( .ip(n1291), .op(n872) );
  nand2_2 U925 ( .ip1(n618), .ip2(n609), .op(n619) );
  nand2_1 U926 ( .ip1(n1526), .ip2(n721), .op(n1487) );
  and2_1 U927 ( .ip1(n1547), .ip2(n1546), .op(n621) );
  nor2_2 U928 ( .ip1(n671), .ip2(n1039), .op(n968) );
  inv_2 U929 ( .ip(n887), .op(n1844) );
  nor2_1 U930 ( .ip1(n1146), .ip2(n1152), .op(n1147) );
  nand2_1 U931 ( .ip1(n1145), .ip2(n1144), .op(n1152) );
  nand2_1 U932 ( .ip1(n1618), .ip2(n1559), .op(n877) );
  nand2_1 U933 ( .ip1(n1618), .ip2(n1617), .op(n1639) );
  nand2_1 U934 ( .ip1(n1143), .ip2(n1612), .op(n1144) );
  nand2_2 U935 ( .ip1(n691), .ip2(n690), .op(n622) );
  nand2_2 U936 ( .ip1(n691), .ip2(n690), .op(n623) );
  nand2_2 U937 ( .ip1(n691), .ip2(n690), .op(n1852) );
  nand2_2 U938 ( .ip1(n685), .ip2(n1833), .op(n691) );
  inv_1 U939 ( .ip(n627), .op(n624) );
  or2_1 U940 ( .ip1(n625), .ip2(n709), .op(n759) );
  nand2_1 U941 ( .ip1(n566), .ip2(n799), .op(n627) );
  inv_1 U942 ( .ip(n1128), .op(n628) );
  inv_1 U943 ( .ip(n611), .op(n855) );
  nand2_1 U944 ( .ip1(n1138), .ip2(n1137), .op(n1558) );
  inv_1 U945 ( .ip(n1655), .op(n629) );
  inv_1 U946 ( .ip(n1667), .op(n630) );
  inv_1 U947 ( .ip(n878), .op(n879) );
  nand2_1 U948 ( .ip1(n876), .ip2(n877), .op(n878) );
  nor2_1 U949 ( .ip1(n775), .ip2(n774), .op(n631) );
  nor2_1 U950 ( .ip1(n1486), .ip2(n773), .op(n632) );
  nor2_1 U951 ( .ip1(n1486), .ip2(n597), .op(n780) );
  nand2_1 U952 ( .ip1(n858), .ip2(partialQ[10]), .op(n633) );
  nand2_1 U953 ( .ip1(n858), .ip2(partialQ[10]), .op(n1599) );
  nand2_2 U954 ( .ip1(counter2Q[3]), .ip2(counter2Q[6]), .op(n677) );
  nand2_1 U955 ( .ip1(n792), .ip2(n793), .op(n798) );
  nand2_1 U956 ( .ip1(n1594), .ip2(n859), .op(n634) );
  nand2_1 U957 ( .ip1(n1594), .ip2(n859), .op(n856) );
  nand2_1 U958 ( .ip1(n879), .ip2(n880), .op(n884) );
  inv_1 U959 ( .ip(n1292), .op(n635) );
  nand2_1 U960 ( .ip1(n568), .ip2(n741), .op(n738) );
  inv_1 U961 ( .ip(n1131), .op(n636) );
  nand2_4 U962 ( .ip1(n1527), .ip2(n1272), .op(n774) );
  nand2_2 U963 ( .ip1(n785), .ip2(n786), .op(n1527) );
  nand2_1 U964 ( .ip1(n802), .ip2(n862), .op(n864) );
  nand2_2 U965 ( .ip1(n628), .ip2(n613), .op(n637) );
  nand2_1 U966 ( .ip1(n613), .ip2(n855), .op(n1142) );
  or2_1 U967 ( .ip1(n636), .ip2(n638), .op(n1265) );
  inv_1 U968 ( .ip(n840), .op(n640) );
  nand2_2 U969 ( .ip1(n733), .ip2(result2[3]), .op(n727) );
  inv_1 U970 ( .ip(n738), .op(n1815) );
  nor2_2 U971 ( .ip1(n1624), .ip2(n716), .op(n777) );
  inv_1 U972 ( .ip(n1624), .op(n1131) );
  inv_2 U973 ( .ip(n620), .op(n840) );
  or2_1 U974 ( .ip1(n810), .ip2(n620), .op(n641) );
  inv_2 U975 ( .ip(n641), .op(n1292) );
  inv_4 U976 ( .ip(n642), .op(n1832) );
  inv_1 U977 ( .ip(n807), .op(n804) );
  nand2_2 U978 ( .ip1(n802), .ip2(n803), .op(n807) );
  nand2_1 U979 ( .ip1(n1262), .ip2(n863), .op(n1263) );
  nand2_2 U980 ( .ip1(n807), .ip2(n806), .op(n1549) );
  xnor2_2 U981 ( .ip1(n643), .ip2(n1525), .op(n1274) );
  or2_1 U982 ( .ip1(n1535), .ip2(n1273), .op(n643) );
  inv_4 U983 ( .ip(n739), .op(n1162) );
  inv_1 U984 ( .ip(n647), .op(n644) );
  inv_2 U985 ( .ip(n769), .op(n1297) );
  nand2_2 U986 ( .ip1(n743), .ip2(n744), .op(n769) );
  nand2_1 U987 ( .ip1(n644), .ip2(n735), .op(n1791) );
  nor2_2 U988 ( .ip1(counter2Q[14]), .ip2(counter2Q[15]), .op(n646) );
  nor2_2 U989 ( .ip1(counter2Q[15]), .ip2(counter2Q[14]), .op(n700) );
  inv_1 U990 ( .ip(n736), .op(n647) );
  buf_4 U991 ( .ip(n733), .op(n725) );
  nand2_4 U992 ( .ip1(n725), .ip2(result2[2]), .op(n739) );
  nor2_4 U993 ( .ip1(n851), .ip2(n706), .op(n707) );
  nor2_2 U994 ( .ip1(counter2Q[8]), .ip2(counter2Q[4]), .op(n699) );
  nor2_1 U995 ( .ip1(n620), .ip2(n838), .op(n685) );
  nor2_4 U996 ( .ip1(counter2Q[0]), .ip2(counter2Q[12]), .op(n679) );
  nand2_1 U997 ( .ip1(n896), .ip2(n1844), .op(n897) );
  inv_1 U998 ( .ip(n1866), .op(n896) );
  inv_1 U999 ( .ip(n990), .op(n992) );
  or2_1 U1000 ( .ip1(n996), .ip2(n1659), .op(n991) );
  nor2_1 U1001 ( .ip1(n1707), .ip2(n1712), .op(n997) );
  nand2_1 U1002 ( .ip1(doB[8]), .ip2(n1880), .op(n1841) );
  nand2_1 U1003 ( .ip1(n768), .ip2(n763), .op(n772) );
  inv_1 U1004 ( .ip(n899), .op(n900) );
  and2_1 U1005 ( .ip1(doB[14]), .ip2(n1844), .op(n1843) );
  nand3_1 U1006 ( .ip1(\mult/counterQ [3]), .ip2(n1864), .ip3(n1863), .op(
        n1839) );
  nand2_1 U1007 ( .ip1(partialQ[13]), .ip2(n842), .op(n1139) );
  inv_2 U1008 ( .ip(n800), .op(n1622) );
  inv_1 U1009 ( .ip(n847), .op(n849) );
  inv_1 U1010 ( .ip(n1468), .op(n1319) );
  nand2_1 U1011 ( .ip1(n669), .ip2(n1535), .op(n721) );
  nand2_1 U1012 ( .ip1(n661), .ip2(n1638), .op(n1627) );
  mux2_1 U1013 ( .ip1(doA[15]), .ip2(doA[14]), .s(n1853), .op(n1897) );
  nand2_1 U1014 ( .ip1(n997), .ip2(n1708), .op(n1765) );
  nand2_2 U1015 ( .ip1(n936), .ip2(n935), .op(n999) );
  inv_1 U1016 ( .ip(n906), .op(n908) );
  inv_1 U1017 ( .ip(n1036), .op(n975) );
  mux2_1 U1018 ( .ip1(doA[13]), .ip2(doA[12]), .s(n1853), .op(n1894) );
  mux2_1 U1019 ( .ip1(doA[11]), .ip2(doA[10]), .s(n1853), .op(n1891) );
  nand2_1 U1020 ( .ip1(n957), .ip2(n956), .op(n958) );
  nand2_2 U1021 ( .ip1(n566), .ip2(n799), .op(n1291) );
  inv_1 U1022 ( .ip(aAQ[0]), .op(n1924) );
  nand2_1 U1023 ( .ip1(n646), .ip2(n699), .op(n704) );
  nand2_1 U1024 ( .ip1(n1140), .ip2(n1139), .op(n1620) );
  inv_1 U1025 ( .ip(n1088), .op(n1091) );
  nand2_1 U1026 ( .ip1(n788), .ip2(n787), .op(n793) );
  nand2_1 U1027 ( .ip1(n791), .ip2(n669), .op(n792) );
  and2_1 U1028 ( .ip1(\mult/storeQ [9]), .ip2(\mult/productQ [9]), .op(n990)
         );
  nor2_2 U1029 ( .ip1(\mult/productQ [9]), .ip2(\mult/storeQ [9]), .op(n996)
         );
  nand2_1 U1030 ( .ip1(n1619), .ip2(n1620), .op(n1637) );
  nand2_1 U1031 ( .ip1(n1626), .ip2(n1625), .op(n1633) );
  inv_1 U1032 ( .ip(n1695), .op(n931) );
  inv_1 U1033 ( .ip(n1374), .op(n1777) );
  mux2_1 U1034 ( .ip1(doA[12]), .ip2(doA[11]), .s(n1853), .op(n1893) );
  mux2_1 U1035 ( .ip1(doA[14]), .ip2(doA[13]), .s(n1853), .op(n1896) );
  mux2_1 U1036 ( .ip1(doA[10]), .ip2(doA[9]), .s(n1853), .op(n1890) );
  mux2_1 U1037 ( .ip1(doA[9]), .ip2(doA[8]), .s(n1853), .op(n1889) );
  nand2_1 U1038 ( .ip1(n726), .ip2(n1163), .op(n1819) );
  inv_1 U1039 ( .ip(n1161), .op(n1821) );
  inv_1 U1040 ( .ip(n1484), .op(n722) );
  inv_1 U1041 ( .ip(n1693), .op(n1694) );
  xnor2_1 U1042 ( .ip1(n1061), .ip2(n1060), .op(n1062) );
  nand2_2 U1043 ( .ip1(n1185), .ip2(n1184), .op(n1681) );
  inv_1 U1044 ( .ip(n825), .op(n826) );
  inv_1 U1045 ( .ip(n945), .op(n946) );
  and2_1 U1046 ( .ip1(aAQ[1]), .ip2(aAQ[0]), .op(n1926) );
  or2_1 U1047 ( .ip1(n1108), .ip2(n1078), .op(n1082) );
  xnor2_1 U1048 ( .ip1(n1771), .ip2(n1770), .op(n1772) );
  nand2_1 U1049 ( .ip1(n903), .ip2(n906), .op(n912) );
  nand2_1 U1050 ( .ip1(n965), .ip2(n667), .op(n973) );
  nand2_1 U1051 ( .ip1(n1384), .ip2(\mult/counterQ [3]), .op(n965) );
  nand3_1 U1052 ( .ip1(n963), .ip2(n962), .ip3(n961), .op(n964) );
  nor2_1 U1053 ( .ip1(n1601), .ip2(n1600), .op(n1602) );
  mux2_1 U1054 ( .ip1(n1190), .ip2(n1237), .s(n671), .op(n526) );
  nor2_1 U1055 ( .ip1(n838), .ip2(n837), .op(n839) );
  inv_1 U1056 ( .ip(doB[2]), .op(n1871) );
  and2_1 U1057 ( .ip1(n733), .ip2(result2[6]), .op(n718) );
  inv_1 U1058 ( .ip(n752), .op(n778) );
  inv_1 U1059 ( .ip(n785), .op(n788) );
  nand2_1 U1060 ( .ip1(result2[15]), .ip2(n1622), .op(n1623) );
  inv_1 U1061 ( .ip(n928), .op(n932) );
  nor2_1 U1062 ( .ip1(n1635), .ip2(n873), .op(n874) );
  nand2_1 U1063 ( .ip1(n873), .ip2(n1833), .op(n865) );
  nand2_1 U1064 ( .ip1(n720), .ip2(n746), .op(n790) );
  inv_1 U1065 ( .ip(n1522), .op(n720) );
  inv_1 U1066 ( .ip(n1526), .op(n1529) );
  nand2_1 U1067 ( .ip1(n1525), .ip2(n1524), .op(n1534) );
  nand2_1 U1068 ( .ip1(n1559), .ip2(n1558), .op(n1563) );
  and2_1 U1069 ( .ip1(n1638), .ip2(n1637), .op(n1640) );
  inv_1 U1070 ( .ip(doA[0]), .op(n1874) );
  nor2_1 U1071 ( .ip1(n1313), .ip2(n1312), .op(n1347) );
  inv_1 U1072 ( .ip(n1499), .op(n1711) );
  nand2_1 U1073 ( .ip1(n985), .ip2(n984), .op(n995) );
  nor2_1 U1074 ( .ip1(n1743), .ip2(n983), .op(n984) );
  and2_1 U1075 ( .ip1(aBQ[1]), .ip2(aBQ[0]), .op(n1914) );
  inv_1 U1076 ( .ip(n1086), .op(n1087) );
  nor2_1 U1077 ( .ip1(n1086), .ip2(n1012), .op(n1014) );
  nor2_1 U1078 ( .ip1(n1089), .ip2(n1094), .op(n1015) );
  and2_1 U1079 ( .ip1(n1112), .ip2(n1111), .op(n1117) );
  mux2_1 U1080 ( .ip1(doA[8]), .ip2(doA[7]), .s(n1854), .op(n1888) );
  nand2_1 U1081 ( .ip1(n1034), .ip2(n1512), .op(n1040) );
  inv_1 U1082 ( .ip(n1487), .op(n1492) );
  nor2_2 U1083 ( .ip1(n780), .ip2(n1484), .op(n1493) );
  inv_1 U1084 ( .ip(n808), .op(n809) );
  nor2_1 U1085 ( .ip1(n653), .ip2(n813), .op(n817) );
  or2_1 U1086 ( .ip1(n1292), .ip2(n1635), .op(n813) );
  inv_1 U1087 ( .ip(n870), .op(n882) );
  inv_1 U1088 ( .ip(n1534), .op(n1531) );
  nor2_2 U1089 ( .ip1(n789), .ip2(n790), .op(n1535) );
  nor2_1 U1090 ( .ip1(n1560), .ip2(n1567), .op(n1561) );
  or2_1 U1091 ( .ip1(n1563), .ip2(n1635), .op(n1560) );
  nand2_1 U1092 ( .ip1(n1175), .ip2(\mult/counterQ [1]), .op(n887) );
  nand2_1 U1093 ( .ip1(n1825), .ip2(partialQ[14]), .op(n1153) );
  inv_1 U1094 ( .ip(n1637), .op(n1628) );
  nor2_1 U1095 ( .ip1(n1661), .ip2(n1660), .op(n1662) );
  nor2_1 U1096 ( .ip1(n1707), .ip2(n1706), .op(n1718) );
  nor2_1 U1097 ( .ip1(n1712), .ip2(n1714), .op(n1502) );
  inv_1 U1098 ( .ip(aBQ[0]), .op(n1915) );
  inv_1 U1099 ( .ip(n820), .op(n821) );
  inv_1 U1100 ( .ip(aAQ[6]), .op(n1944) );
  inv_1 U1101 ( .ip(n831), .op(n832) );
  inv_1 U1102 ( .ip(aBQ[6]), .op(n1902) );
  or2_1 U1103 ( .ip1(n1099), .ip2(n1100), .op(n1104) );
  or2_1 U1104 ( .ip1(n1014), .ip2(n1015), .op(n1017) );
  or2_1 U1105 ( .ip1(n1116), .ip2(n1117), .op(n1121) );
  nor2_1 U1106 ( .ip1(n1754), .ip2(n1753), .op(n1755) );
  nor2_1 U1107 ( .ip1(n1744), .ip2(n1743), .op(n1758) );
  nor2_1 U1108 ( .ip1(n1749), .ip2(n1736), .op(n1737) );
  nand2_1 U1109 ( .ip1(n1373), .ip2(n1372), .op(n1378) );
  nand2_1 U1110 ( .ip1(n1370), .ip2(n1369), .op(n1380) );
  nor2_1 U1111 ( .ip1(n1778), .ip2(n1777), .op(n1782) );
  nand4_1 U1112 ( .ip1(n1474), .ip2(n1473), .ip3(n1472), .ip4(n1471), .op(
        n1475) );
  nor2_1 U1113 ( .ip1(n1447), .ip2(n1446), .op(n1448) );
  nand3_1 U1114 ( .ip1(n1459), .ip2(n1458), .ip3(n1457), .op(n1460) );
  inv_1 U1115 ( .ip(reset), .op(n1181) );
  nand2_1 U1116 ( .ip1(n1822), .ip2(n1161), .op(n1823) );
  nand2_1 U1117 ( .ip1(n1525), .ip2(n1483), .op(n1495) );
  inv_1 U1118 ( .ip(n596), .op(n1483) );
  inv_1 U1119 ( .ip(n1495), .op(n1485) );
  nand2_1 U1120 ( .ip1(n724), .ip2(n753), .op(n751) );
  or2_1 U1121 ( .ip1(n763), .ip2(n1295), .op(n1296) );
  inv_1 U1122 ( .ip(n627), .op(n1301) );
  mux2_1 U1123 ( .ip1(n1239), .ip2(n1180), .s(\mult/counterQ [3]), .op(n525)
         );
  xnor2_1 U1124 ( .ip1(n1220), .ip2(n1218), .op(n1219) );
  xnor2_1 U1125 ( .ip1(n1212), .ip2(n1211), .op(n1213) );
  xnor2_1 U1126 ( .ip1(n1223), .ip2(n1222), .op(n1224) );
  xnor2_1 U1127 ( .ip1(n1676), .ip2(n1675), .op(n1677) );
  mux2_1 U1128 ( .ip1(n1386), .ip2(n1385), .s(n1512), .op(n1387) );
  xnor2_1 U1129 ( .ip1(n1684), .ip2(n1683), .op(n1685) );
  nand2_1 U1130 ( .ip1(n1783), .ip2(n1702), .op(n1703) );
  xnor2_1 U1131 ( .ip1(n1653), .ip2(n1652), .op(n1654) );
  nor2_1 U1132 ( .ip1(n1668), .ip2(n1651), .op(n1652) );
  xnor2_1 U1133 ( .ip1(n1657), .ip2(n1656), .op(n1658) );
  nor2_1 U1134 ( .ip1(n1681), .ip2(n1655), .op(n1656) );
  xnor2_1 U1135 ( .ip1(n1670), .ip2(n1669), .op(n1671) );
  nor2_1 U1136 ( .ip1(n1668), .ip2(n1667), .op(n1669) );
  xnor2_1 U1137 ( .ip1(n571), .ip2(n1227), .op(n1228) );
  xnor2_1 U1138 ( .ip1(n1204), .ip2(n1203), .op(n1205) );
  inv_1 U1139 ( .ip(n1235), .op(n1236) );
  inv_1 U1140 ( .ip(n1062), .op(n1063) );
  nand2_1 U1141 ( .ip1(n1075), .ip2(n1074), .op(n489) );
  nand2_1 U1142 ( .ip1(n1070), .ip2(n1069), .op(n488) );
  nand2_1 U1143 ( .ip1(n1783), .ip2(n538), .op(n1070) );
  xnor2_1 U1144 ( .ip1(n1207), .ip2(n1206), .op(n1208) );
  nand2_1 U1145 ( .ip1(n948), .ip2(n947), .op(n1931) );
  inv_1 U1146 ( .ip(n1248), .op(n1249) );
  nor2_1 U1147 ( .ip1(n1171), .ip2(n1170), .op(n1957) );
  nand2_1 U1148 ( .ip1(n1760), .ip2(\mult/productQ [20]), .op(n1084) );
  inv_1 U1149 ( .ip(n1772), .op(n1773) );
  nand3_1 U1150 ( .ip1(n1283), .ip2(n671), .ip3(n1418), .op(n1290) );
  nand2_1 U1151 ( .ip1(n978), .ip2(n1518), .op(n979) );
  nor2_1 U1152 ( .ip1(n973), .ip2(n972), .op(n978) );
  inv_1 U1153 ( .ip(n1126), .op(N318) );
  nor2_1 U1154 ( .ip1(n588), .ip2(n1635), .op(n1125) );
  inv_2 U1155 ( .ip(n733), .op(n800) );
  and2_1 U1156 ( .ip1(n1135), .ip2(n653), .op(n650) );
  or2_1 U1157 ( .ip1(partialQ[13]), .ip2(result2[13]), .op(n654) );
  and2_4 U1158 ( .ip1(\mult/counterQ [3]), .ip2(n1506), .op(n655) );
  nand2_1 U1159 ( .ip1(\mult/counterQ [2]), .ip2(\mult/counterQ [3]), .op(n656) );
  and2_1 U1160 ( .ip1(n812), .ip2(n811), .op(n657) );
  and2_1 U1161 ( .ip1(n768), .ip2(n1296), .op(n659) );
  and2_1 U1162 ( .ip1(n1552), .ip2(n1833), .op(n660) );
  nand2_1 U1163 ( .ip1(doB[10]), .ip2(n1844), .op(n662) );
  and2_1 U1164 ( .ip1(n1037), .ip2(n1036), .op(n663) );
  and2_1 U1165 ( .ip1(n1422), .ip2(\mult/counterQ [3]), .op(n664) );
  and2_1 U1166 ( .ip1(n1789), .ip2(n734), .op(n665) );
  and2_1 U1167 ( .ip1(n1634), .ip2(n1633), .op(n666) );
  or2_1 U1168 ( .ip1(n539), .ip2(n964), .op(n667) );
  and2_1 U1169 ( .ip1(n1137), .ip2(n654), .op(n668) );
  nand2_2 U1170 ( .ip1(n759), .ip2(n1304), .op(n1548) );
  or2_1 U1171 ( .ip1(partialQ[5]), .ip2(result2[5]), .op(n669) );
  inv_1 U1172 ( .ip(partialQ[13]), .op(n1136) );
  inv_1 U1173 ( .ip(n1371), .op(n1779) );
  and2_1 U1174 ( .ip1(n1195), .ip2(n1192), .op(n670) );
  nand2_1 U1176 ( .ip1(n673), .ip2(n672), .op(n676) );
  nor2_2 U1177 ( .ip1(counter2Q[10]), .ip2(counter2Q[5]), .op(n701) );
  nand2_1 U1178 ( .ip1(n701), .ip2(n674), .op(n675) );
  nor2_2 U1179 ( .ip1(n675), .ip2(n676), .op(n853) );
  inv_2 U1180 ( .ip(n677), .op(n702) );
  nand2_2 U1181 ( .ip1(n700), .ip2(n702), .op(n850) );
  inv_2 U1182 ( .ip(n678), .op(n680) );
  nand2_4 U1183 ( .ip1(n679), .ip2(n680), .op(n851) );
  nand2_4 U1184 ( .ip1(counterQ[3]), .ip2(n683), .op(n733) );
  inv_2 U1185 ( .ip(n733), .op(n838) );
  inv_2 U1186 ( .ip(state[1]), .op(n1586) );
  inv_1 U1187 ( .ip(wrAddr[1]), .op(n695) );
  nand2_1 U1188 ( .ip1(wrAddr[0]), .ip2(n695), .op(n686) );
  nor2_1 U1189 ( .ip1(n686), .ip2(state[1]), .op(n692) );
  or2_1 U1190 ( .ip1(wrAddr[3]), .ip2(wrAddr[2]), .op(n694) );
  nor2_1 U1191 ( .ip1(n694), .ip2(state[0]), .op(n687) );
  nand2_1 U1192 ( .ip1(n692), .ip2(n687), .op(n441) );
  nand2_1 U1193 ( .ip1(n1898), .ip2(n1181), .op(n688) );
  nand2_1 U1194 ( .ip1(n1942), .ip2(n1941), .op(n1270) );
  nand2_1 U1195 ( .ip1(n622), .ip2(n1270), .op(n715) );
  inv_1 U1196 ( .ip(n692), .op(n693) );
  nor2_1 U1197 ( .ip1(n694), .ip2(n693), .op(n698) );
  inv_1 U1198 ( .ip(state[0]), .op(n1169) );
  or4_1 U1199 ( .ip1(wrAddr[3]), .ip2(wrAddr[0]), .ip3(wrAddr[2]), .ip4(n695), 
        .op(n696) );
  nand2_1 U1200 ( .ip1(n1169), .ip2(n696), .op(n697) );
  nand2_1 U1201 ( .ip1(n697), .ip2(n1586), .op(n1170) );
  nand2_2 U1202 ( .ip1(n1170), .ip2(n1181), .op(n1593) );
  or2_1 U1203 ( .ip1(n698), .ip2(n1593), .op(n713) );
  nand2_1 U1204 ( .ip1(n701), .ip2(n702), .op(n703) );
  nor2_2 U1205 ( .ip1(n704), .ip2(n703), .op(n708) );
  nor2_2 U1206 ( .ip1(counter2Q[11]), .ip2(counter2Q[7]), .op(n705) );
  nand2_1 U1207 ( .ip1(n802), .ip2(n1622), .op(n709) );
  inv_4 U1208 ( .ip(n711), .op(n1635) );
  nand2_4 U1209 ( .ip1(n713), .ip2(n712), .op(n714) );
  inv_4 U1210 ( .ip(n714), .op(n1544) );
  nand2_2 U1211 ( .ip1(n715), .ip2(n1544), .op(n1946) );
  inv_1 U1212 ( .ip(partialQ[7]), .op(n752) );
  nand2_1 U1213 ( .ip1(n777), .ip2(partialQ[7]), .op(n781) );
  nand2_1 U1214 ( .ip1(n794), .ip2(n781), .op(n717) );
  nand2_1 U1215 ( .ip1(n717), .ip2(n1833), .op(n754) );
  nor2_1 U1216 ( .ip1(n1635), .ip2(n717), .op(n724) );
  and2_1 U1217 ( .ip1(n1486), .ip2(n597), .op(n1484) );
  nor2_4 U1218 ( .ip1(n838), .ip2(n719), .op(n783) );
  inv_1 U1219 ( .ip(partialQ[5]), .op(n786) );
  inv_1 U1220 ( .ip(n620), .op(n784) );
  nand3_1 U1221 ( .ip1(n840), .ip2(partialQ[5]), .ip3(n783), .op(n1526) );
  inv_1 U1222 ( .ip(partialQ[4]), .op(n1522) );
  inv_2 U1223 ( .ip(result2[4]), .op(n1523) );
  nor2_2 U1224 ( .ip1(n780), .ip2(n723), .op(n753) );
  inv_1 U1225 ( .ip(partialQ[3]), .op(n1814) );
  inv_2 U1226 ( .ip(result2[0]), .op(n765) );
  nand2_2 U1227 ( .ip1(n588), .ip2(n731), .op(n1261) );
  nor2_2 U1228 ( .ip1(n838), .ip2(n734), .op(n762) );
  nand2_2 U1229 ( .ip1(n737), .ip2(n645), .op(n1820) );
  nand2_2 U1230 ( .ip1(n768), .ip2(n1820), .op(n745) );
  nand2_2 U1231 ( .ip1(partialQ[2]), .ip2(n1162), .op(n740) );
  inv_2 U1232 ( .ip(n740), .op(n1160) );
  nand2_2 U1233 ( .ip1(n745), .ip2(n770), .op(n1525) );
  nor2_1 U1234 ( .ip1(partialQ[6]), .ip2(result2[6]), .op(n748) );
  nand2_1 U1235 ( .ip1(n802), .ip2(n746), .op(n747) );
  mux2_1 U1236 ( .ip1(n754), .ip2(n751), .s(n750), .op(n758) );
  nor2_1 U1237 ( .ip1(n752), .ip2(n1593), .op(n756) );
  nor2_1 U1238 ( .ip1(n754), .ip2(n753), .op(n755) );
  nor2_1 U1239 ( .ip1(n756), .ip2(n755), .op(n757) );
  nand2_1 U1240 ( .ip1(n757), .ip2(n758), .op(n450) );
  inv_1 U1241 ( .ip(partialQ[8]), .op(n1304) );
  inv_1 U1242 ( .ip(n1548), .op(n760) );
  inv_2 U1243 ( .ip(n760), .op(n815) );
  nand3_1 U1244 ( .ip1(n735), .ip2(n1131), .ip3(n762), .op(n1294) );
  inv_1 U1245 ( .ip(n1294), .op(n763) );
  nor2_1 U1246 ( .ip1(partialQ[1]), .ip2(result2[1]), .op(n764) );
  inv_1 U1247 ( .ip(n769), .op(n770) );
  nand3_2 U1248 ( .ip1(n771), .ip2(n772), .ip3(n1297), .op(n776) );
  nand2_2 U1249 ( .ip1(n794), .ip2(n795), .op(n775) );
  nor2_4 U1250 ( .ip1(n775), .ip2(n774), .op(n1293) );
  or2_1 U1251 ( .ip1(n778), .ip2(n777), .op(n779) );
  nand2_1 U1252 ( .ip1(n632), .ip2(n779), .op(n782) );
  nand2_2 U1253 ( .ip1(n798), .ip2(n797), .op(n799) );
  nand2_1 U1254 ( .ip1(n609), .ip2(n872), .op(n814) );
  nand3_1 U1255 ( .ip1(n814), .ip2(n815), .ip3(n650), .op(n819) );
  nand2_1 U1256 ( .ip1(result2[8]), .ip2(partialQ[8]), .op(n808) );
  nand2_1 U1257 ( .ip1(n809), .ip2(n733), .op(n810) );
  nand3_1 U1258 ( .ip1(n1292), .ip2(n653), .ip3(n1833), .op(n812) );
  inv_2 U1259 ( .ip(n1593), .op(n1825) );
  nand2_1 U1260 ( .ip1(n1825), .ip2(partialQ[9]), .op(n811) );
  nand2_1 U1261 ( .ip1(n814), .ip2(n815), .op(n816) );
  nand2_1 U1262 ( .ip1(n817), .ip2(n816), .op(n818) );
  nand3_1 U1263 ( .ip1(n818), .ip2(n657), .ip3(n819), .op(n448) );
  nand2_1 U1264 ( .ip1(n622), .ip2(n1950), .op(n820) );
  nor2_1 U1265 ( .ip1(n1946), .ip2(n821), .op(n823) );
  inv_1 U1266 ( .ip(n1947), .op(n822) );
  nand2_1 U1267 ( .ip1(n823), .ip2(n822), .op(n1951) );
  nand2_1 U1268 ( .ip1(n1852), .ip2(n1915), .op(n824) );
  nand2_1 U1269 ( .ip1(n622), .ip2(n1917), .op(n825) );
  nor2_1 U1270 ( .ip1(n1922), .ip2(n826), .op(n828) );
  inv_1 U1271 ( .ip(n1916), .op(n827) );
  nand2_1 U1272 ( .ip1(n828), .ip2(n827), .op(n1918) );
  nor2_1 U1273 ( .ip1(n1917), .ip2(n1900), .op(n829) );
  and2_1 U1274 ( .ip1(n1914), .ip2(n829), .op(n1907) );
  nand2_1 U1275 ( .ip1(n1907), .ip2(n1901), .op(n1268) );
  nand2_1 U1276 ( .ip1(n623), .ip2(n1954), .op(n831) );
  nor2_1 U1277 ( .ip1(n1905), .ip2(n832), .op(n834) );
  inv_1 U1278 ( .ip(n1903), .op(n833) );
  nand2_1 U1279 ( .ip1(n834), .ip2(n833), .op(n1955) );
  nand2_1 U1280 ( .ip1(n1825), .ip2(partialQ[13]), .op(n835) );
  and2_1 U1281 ( .ip1(result2[12]), .ip2(partialQ[12]), .op(n1137) );
  inv_1 U1282 ( .ip(n1558), .op(n843) );
  inv_1 U1283 ( .ip(result2[13]), .op(n837) );
  nand2_1 U1284 ( .ip1(n1159), .ip2(n839), .op(n841) );
  nand2_1 U1285 ( .ip1(n1136), .ip2(n841), .op(n1127) );
  inv_1 U1286 ( .ip(n841), .op(n842) );
  nand2_1 U1287 ( .ip1(n1127), .ip2(n1139), .op(n873) );
  nand2_1 U1288 ( .ip1(n843), .ip2(n881), .op(n844) );
  nand2_1 U1289 ( .ip1(n835), .ip2(n844), .op(n867) );
  nand2_1 U1290 ( .ip1(n588), .ip2(result2[11]), .op(n847) );
  inv_1 U1291 ( .ip(partialQ[10]), .op(n854) );
  nand2_1 U1292 ( .ip1(n857), .ip2(n854), .op(n1587) );
  inv_1 U1293 ( .ip(n857), .op(n858) );
  nor2_2 U1294 ( .ip1(n1591), .ip2(n1599), .op(n860) );
  nor2_1 U1295 ( .ip1(n859), .ip2(n1594), .op(n1590) );
  nor2_2 U1296 ( .ip1(n860), .ip2(n1590), .op(n1141) );
  nand2_2 U1297 ( .ip1(n1141), .ip2(n637), .op(n1618) );
  inv_1 U1298 ( .ip(partialQ[12]), .op(n1566) );
  nand2_2 U1299 ( .ip1(n1566), .ip2(n864), .op(n1559) );
  nor2_1 U1300 ( .ip1(n877), .ip2(n865), .op(n866) );
  nor2_1 U1301 ( .ip1(n867), .ip2(n866), .op(n885) );
  inv_1 U1302 ( .ip(n1559), .op(n868) );
  nand2_1 U1303 ( .ip1(n869), .ip2(n815), .op(n870) );
  nand2_1 U1304 ( .ip1(n874), .ip2(n1558), .op(n875) );
  inv_1 U1305 ( .ip(n875), .op(n876) );
  nand3_1 U1306 ( .ip1(n626), .ip2(n882), .ip3(n881), .op(n883) );
  nand3_1 U1307 ( .ip1(n884), .ip2(n885), .ip3(n883), .op(n444) );
  nand2_1 U1308 ( .ip1(n1892), .ip2(\mult/counterQ [3]), .op(n886) );
  nand2_1 U1309 ( .ip1(n886), .ip2(n1842), .op(n891) );
  inv_4 U1310 ( .ip(\mult/counterQ [0]), .op(n1175) );
  nor2_1 U1311 ( .ip1(n1871), .ip2(\mult/counterQ [2]), .op(n888) );
  nand2_1 U1312 ( .ip1(n1844), .ip2(n888), .op(n889) );
  nand2_1 U1313 ( .ip1(n1872), .ip2(n889), .op(n890) );
  nor2_2 U1314 ( .ip1(n891), .ip2(n890), .op(n892) );
  nand3_2 U1315 ( .ip1(n649), .ip2(n662), .ip3(n1841), .op(n967) );
  nand2_1 U1316 ( .ip1(n907), .ip2(n967), .op(n950) );
  buf_1 U1317 ( .ip(\mult/counterQ [1]), .op(n893) );
  nor2_2 U1318 ( .ip1(n1867), .ip2(n1443), .op(n895) );
  inv_1 U1319 ( .ip(n1846), .op(n894) );
  inv_1 U1320 ( .ip(n1870), .op(n1198) );
  nor2_1 U1321 ( .ip1(n1865), .ip2(n1198), .op(n899) );
  inv_2 U1322 ( .ip(\mult/counterQ [5]), .op(n1195) );
  nand2_2 U1323 ( .ip1(\mult/state [0]), .ip2(n1181), .op(n951) );
  inv_2 U1324 ( .ip(n951), .op(n1192) );
  nand3_2 U1325 ( .ip1(n950), .ip2(n949), .ip3(n670), .op(n905) );
  and2_2 U1326 ( .ip1(\mult/state [1]), .ip2(n1181), .op(n952) );
  inv_1 U1327 ( .ip(n952), .op(n904) );
  nand2_4 U1328 ( .ip1(n905), .ip2(n904), .op(n1760) );
  nand2_1 U1329 ( .ip1(n1760), .ip2(\mult/productQ [9]), .op(n943) );
  nor2_1 U1330 ( .ip1(n951), .ip2(n952), .op(n906) );
  nand3_1 U1331 ( .ip1(n906), .ip2(n1036), .ip3(n595), .op(n913) );
  inv_2 U1332 ( .ip(n907), .op(n1039) );
  nor2_2 U1333 ( .ip1(n908), .ip2(n1039), .op(n910) );
  buf_1 U1334 ( .ip(n967), .op(n909) );
  nand2_2 U1335 ( .ip1(n910), .ip2(n909), .op(n911) );
  nand3_4 U1336 ( .ip1(n913), .ip2(n912), .ip3(n911), .op(n1774) );
  buf_4 U1337 ( .ip(n1774), .op(n1810) );
  nor2_1 U1338 ( .ip1(n996), .ip2(n990), .op(n940) );
  nor2_1 U1339 ( .ip1(\mult/storeQ [2]), .ip2(\mult/productQ [2]), .op(n1363)
         );
  nor2_2 U1340 ( .ip1(\mult/storeQ [3]), .ip2(\mult/productQ [3]), .op(n1057)
         );
  nor2_1 U1341 ( .ip1(n1363), .ip2(n1057), .op(n917) );
  nand2_1 U1342 ( .ip1(\mult/storeQ [1]), .ip2(\mult/productQ [1]), .op(n1066)
         );
  and2_2 U1343 ( .ip1(\mult/storeQ [0]), .ip2(\mult/productQ [0]), .op(n1071)
         );
  nand2_2 U1344 ( .ip1(n915), .ip2(n914), .op(n1067) );
  nand2_2 U1345 ( .ip1(n1071), .ip2(n1067), .op(n916) );
  nand2_2 U1346 ( .ip1(n1066), .ip2(n916), .op(n1364) );
  nand2_2 U1347 ( .ip1(n917), .ip2(n1364), .op(n920) );
  and2_1 U1348 ( .ip1(\mult/productQ [3]), .ip2(\mult/storeQ [3]), .op(n1056)
         );
  nand2_1 U1349 ( .ip1(\mult/productQ [2]), .ip2(\mult/storeQ [2]), .op(n1361)
         );
  nand2_2 U1350 ( .ip1(n920), .ip2(n919), .op(n1697) );
  inv_1 U1351 ( .ip(\mult/productQ [6]), .op(n922) );
  inv_1 U1352 ( .ip(\mult/storeQ [6]), .op(n921) );
  inv_1 U1353 ( .ip(\mult/productQ [7]), .op(n924) );
  inv_1 U1354 ( .ip(\mult/storeQ [7]), .op(n923) );
  nand2_1 U1355 ( .ip1(n1374), .ip2(n1370), .op(n928) );
  or2_1 U1356 ( .ip1(\mult/storeQ [4]), .ip2(\mult/productQ [4]), .op(n1696)
         );
  nand2_1 U1357 ( .ip1(n1696), .ip2(n1693), .op(n1375) );
  nor2_1 U1358 ( .ip1(n928), .ip2(n1375), .op(n925) );
  nand2_2 U1359 ( .ip1(n1697), .ip2(n925), .op(n936) );
  and2_1 U1360 ( .ip1(\mult/storeQ [6]), .ip2(\mult/productQ [6]), .op(n1778)
         );
  nand2_1 U1361 ( .ip1(n1370), .ip2(n1778), .op(n926) );
  nand2_1 U1362 ( .ip1(\mult/storeQ [7]), .ip2(\mult/productQ [7]), .op(n1369)
         );
  and2_1 U1363 ( .ip1(\mult/productQ [5]), .ip2(\mult/storeQ [5]), .op(n1695)
         );
  nor2_2 U1364 ( .ip1(\mult/storeQ [8]), .ip2(\mult/productQ [8]), .op(n1661)
         );
  inv_1 U1365 ( .ip(n1661), .op(n937) );
  nand2_1 U1366 ( .ip1(n1767), .ip2(n937), .op(n938) );
  nand2_1 U1367 ( .ip1(\mult/storeQ [8]), .ip2(\mult/productQ [8]), .op(n1659)
         );
  nand2_1 U1368 ( .ip1(n938), .ip2(n1659), .op(n939) );
  xor2_1 U1369 ( .ip1(n940), .ip2(n939), .op(n941) );
  nand2_4 U1370 ( .ip1(n1783), .ip2(n941), .op(n942) );
  buf_2 U1371 ( .ip(\mult/counterQ [1]), .op(n1851) );
  nor2_1 U1372 ( .ip1(n1947), .ip2(n1946), .op(n1835) );
  nor2_1 U1373 ( .ip1(n1922), .ip2(n1916), .op(n1836) );
  nor2_1 U1374 ( .ip1(n1905), .ip2(n1903), .op(n1837) );
  nand2_1 U1375 ( .ip1(n622), .ip2(n1924), .op(n944) );
  nand2_1 U1376 ( .ip1(n944), .ip2(n1544), .op(n1927) );
  inv_1 U1377 ( .ip(n1927), .op(n948) );
  nand2_1 U1378 ( .ip1(n623), .ip2(n1930), .op(n945) );
  nand3_1 U1379 ( .ip1(n950), .ip2(n949), .ip3(n1192), .op(n953) );
  nor2_2 U1380 ( .ip1(n951), .ip2(n1195), .op(n1191) );
  nor2_2 U1381 ( .ip1(n1191), .ip2(n952), .op(n1174) );
  nand2_2 U1382 ( .ip1(n953), .ip2(n1174), .op(n1022) );
  nand2_1 U1383 ( .ip1(n1480), .ip2(\mult/storeQ [17]), .op(n980) );
  inv_2 U1384 ( .ip(n1175), .op(n1853) );
  nor2_1 U1385 ( .ip1(n1443), .ip2(n1318), .op(n960) );
  buf_1 U1386 ( .ip(n1851), .op(n1349) );
  inv_2 U1387 ( .ip(n1469), .op(n1343) );
  nor2_1 U1388 ( .ip1(n1343), .ip2(n1342), .op(n959) );
  inv_1 U1389 ( .ip(n1406), .op(n954) );
  inv_2 U1390 ( .ip(\mult/counterQ [1]), .op(n1445) );
  buf_2 U1391 ( .ip(n1850), .op(n1468) );
  nand2_1 U1392 ( .ip1(n954), .ip2(n1468), .op(n957) );
  nor2_2 U1393 ( .ip1(n1349), .ip2(\mult/counterQ [2]), .op(n955) );
  nand2_1 U1394 ( .ip1(n1889), .ip2(n1470), .op(n956) );
  nor3_2 U1395 ( .ip1(n960), .ip2(n959), .ip3(n958), .op(n1384) );
  nand2_1 U1396 ( .ip1(n1894), .ip2(n1469), .op(n963) );
  nand2_1 U1397 ( .ip1(n1891), .ip2(n1511), .op(n962) );
  nand2_1 U1398 ( .ip1(n1897), .ip2(n1468), .op(n961) );
  inv_2 U1399 ( .ip(n1470), .op(n1317) );
  nand2_2 U1400 ( .ip1(n1192), .ip2(n1174), .op(n1177) );
  inv_2 U1401 ( .ip(n1177), .op(n966) );
  nand2_2 U1402 ( .ip1(n968), .ip2(n1042), .op(n971) );
  nand2_2 U1403 ( .ip1(n966), .ip2(n1840), .op(n1033) );
  inv_2 U1404 ( .ip(n1033), .op(n969) );
  nand2_2 U1405 ( .ip1(n652), .ip2(n969), .op(n970) );
  nand2_4 U1406 ( .ip1(n971), .ip2(n970), .op(n1506) );
  nor2_1 U1407 ( .ip1(n1386), .ip2(n1506), .op(n972) );
  nor2_1 U1408 ( .ip1(n1039), .ip2(n974), .op(n977) );
  nor2_2 U1409 ( .ip1(n975), .ip2(n1033), .op(n976) );
  nor2_2 U1410 ( .ip1(n977), .ip2(n976), .op(n1030) );
  nor2_2 U1411 ( .ip1(n1030), .ip2(\mult/counterQ [3]), .op(n1283) );
  nand2_1 U1412 ( .ip1(n980), .ip2(n979), .op(n504) );
  inv_4 U1413 ( .ip(n1175), .op(n1854) );
  nor2_2 U1414 ( .ip1(n1854), .ip2(n1851), .op(n1880) );
  nor2_1 U1415 ( .ip1(\mult/storeQ [13]), .ip2(\mult/productQ [13]), .op(n1724) );
  inv_1 U1416 ( .ip(n1724), .op(n981) );
  and2_1 U1417 ( .ip1(\mult/productQ [12]), .ip2(\mult/storeQ [12]), .op(n1763) );
  nand2_1 U1418 ( .ip1(n981), .ip2(n1763), .op(n982) );
  nand2_1 U1419 ( .ip1(\mult/storeQ [13]), .ip2(\mult/productQ [13]), .op(
        n1722) );
  nand2_1 U1420 ( .ip1(n982), .ip2(n1722), .op(n1749) );
  nor2_1 U1421 ( .ip1(\mult/storeQ [14]), .ip2(\mult/productQ [14]), .op(n1745) );
  nor2_1 U1422 ( .ip1(\mult/storeQ [15]), .ip2(\mult/productQ [15]), .op(n1744) );
  nor2_1 U1423 ( .ip1(n1745), .ip2(n1744), .op(n986) );
  nand2_1 U1424 ( .ip1(n1749), .ip2(n986), .op(n985) );
  and2_1 U1425 ( .ip1(\mult/productQ [15]), .ip2(\mult/storeQ [15]), .op(n1743) );
  nand2_1 U1426 ( .ip1(\mult/storeQ [14]), .ip2(\mult/productQ [14]), .op(
        n1750) );
  nor2_1 U1427 ( .ip1(n1750), .ip2(n1744), .op(n983) );
  nor2_1 U1428 ( .ip1(\mult/storeQ [12]), .ip2(\mult/productQ [12]), .op(n1764) );
  nor2_1 U1429 ( .ip1(n1724), .ip2(n1764), .op(n1746) );
  nand2_1 U1430 ( .ip1(n986), .ip2(n1746), .op(n998) );
  nor2_2 U1431 ( .ip1(\mult/storeQ [11]), .ip2(\mult/productQ [11]), .op(n1707) );
  inv_1 U1432 ( .ip(n1707), .op(n987) );
  and2_1 U1433 ( .ip1(\mult/productQ [10]), .ip2(\mult/storeQ [10]), .op(n1714) );
  nand2_1 U1434 ( .ip1(n987), .ip2(n1714), .op(n988) );
  nand2_1 U1435 ( .ip1(\mult/storeQ [11]), .ip2(\mult/productQ [11]), .op(
        n1705) );
  nor2_2 U1436 ( .ip1(\mult/storeQ [10]), .ip2(\mult/productQ [10]), .op(n1712) );
  and2_2 U1437 ( .ip1(n989), .ip2(n993), .op(n1768) );
  nor2_2 U1438 ( .ip1(n998), .ip2(n1768), .op(n994) );
  nor2_1 U1439 ( .ip1(n996), .ip2(n1661), .op(n1708) );
  nor2_1 U1440 ( .ip1(n998), .ip2(n1765), .op(n1000) );
  or2_1 U1441 ( .ip1(\mult/storeQ [20]), .ip2(\mult/productQ [20]), .op(n1076)
         );
  or2_1 U1442 ( .ip1(\mult/storeQ [21]), .ip2(\mult/productQ [21]), .op(n1112)
         );
  nand2_1 U1443 ( .ip1(n1076), .ip2(n1112), .op(n1088) );
  nor2_1 U1444 ( .ip1(\mult/storeQ [16]), .ip2(\mult/productQ [16]), .op(n1688) );
  nor2_1 U1445 ( .ip1(\mult/storeQ [17]), .ip2(\mult/productQ [17]), .op(n1575) );
  nor2_1 U1446 ( .ip1(n1688), .ip2(n1575), .op(n1799) );
  nor2_1 U1447 ( .ip1(\mult/storeQ [18]), .ip2(\mult/productQ [18]), .op(n1804) );
  nor2_1 U1448 ( .ip1(\mult/storeQ [19]), .ip2(\mult/productQ [19]), .op(n1798) );
  nor2_1 U1449 ( .ip1(n1804), .ip2(n1798), .op(n1007) );
  nand2_1 U1450 ( .ip1(n1799), .ip2(n1007), .op(n1113) );
  nor2_1 U1451 ( .ip1(n1088), .ip2(n1113), .op(n1003) );
  nand2_1 U1452 ( .ip1(n1802), .ip2(n1003), .op(n1013) );
  nor2_1 U1453 ( .ip1(\mult/storeQ [22]), .ip2(\mult/productQ [22]), .op(n1089) );
  and2_1 U1454 ( .ip1(\mult/productQ [22]), .ip2(\mult/storeQ [22]), .op(n1094) );
  or2_1 U1455 ( .ip1(n1013), .ip2(n1015), .op(n1018) );
  and2_1 U1456 ( .ip1(\mult/productQ [20]), .ip2(\mult/storeQ [20]), .op(n1110) );
  nand2_1 U1457 ( .ip1(n1112), .ip2(n1110), .op(n1004) );
  nand2_1 U1458 ( .ip1(\mult/productQ [21]), .ip2(\mult/storeQ [21]), .op(
        n1111) );
  nand2_1 U1459 ( .ip1(n1004), .ip2(n1111), .op(n1086) );
  inv_1 U1460 ( .ip(n1798), .op(n1005) );
  and2_1 U1461 ( .ip1(\mult/productQ [18]), .ip2(\mult/storeQ [18]), .op(n1806) );
  nand2_1 U1462 ( .ip1(n1005), .ip2(n1806), .op(n1006) );
  nand2_1 U1463 ( .ip1(\mult/productQ [19]), .ip2(\mult/storeQ [19]), .op(
        n1796) );
  nand2_1 U1464 ( .ip1(n1006), .ip2(n1796), .op(n1011) );
  inv_1 U1465 ( .ip(n1007), .op(n1009) );
  and2_1 U1466 ( .ip1(\mult/productQ [17]), .ip2(\mult/storeQ [17]), .op(n1574) );
  nand2_1 U1467 ( .ip1(\mult/storeQ [16]), .ip2(\mult/productQ [16]), .op(
        n1686) );
  nor2_1 U1468 ( .ip1(n1686), .ip2(n1575), .op(n1008) );
  nor2_2 U1469 ( .ip1(n1011), .ip2(n1010), .op(n1108) );
  nor2_1 U1470 ( .ip1(n1088), .ip2(n1108), .op(n1012) );
  nand3_1 U1471 ( .ip1(n1015), .ip2(n1014), .ip3(n1013), .op(n1016) );
  nand3_1 U1472 ( .ip1(n1018), .ip2(n1017), .ip3(n1016), .op(n1019) );
  nand2_1 U1473 ( .ip1(n1019), .ip2(n573), .op(n1021) );
  nand2_1 U1474 ( .ip1(n1760), .ip2(\mult/productQ [22]), .op(n1020) );
  nand2_1 U1475 ( .ip1(n1021), .ip2(n1020), .op(n467) );
  nand2_1 U1476 ( .ip1(n1519), .ip2(\mult/storeQ [22]), .op(n1055) );
  not_ab_or_c_or_d U1477 ( .ip1(n1445), .ip2(n1883), .ip3(n1882), .ip4(n1892), 
        .op(n1028) );
  inv_1 U1478 ( .ip(n1886), .op(n1023) );
  nand2_1 U1479 ( .ip1(n1023), .ip2(n1468), .op(n1026) );
  inv_1 U1480 ( .ip(n1887), .op(n1024) );
  nand2_1 U1481 ( .ip1(n1024), .ip2(n1470), .op(n1025) );
  nand2_1 U1482 ( .ip1(n1026), .ip2(n1025), .op(n1027) );
  and2_1 U1483 ( .ip1(n1895), .ip2(n1851), .op(n1456) );
  nand2_1 U1484 ( .ip1(n1456), .ip2(\mult/counterQ [2]), .op(n1029) );
  nand2_1 U1485 ( .ip1(n1029), .ip2(n1034), .op(n1045) );
  nand2_1 U1486 ( .ip1(n651), .ip2(n1512), .op(n1031) );
  or2_1 U1487 ( .ip1(n1031), .ip2(n1030), .op(n1032) );
  inv_1 U1488 ( .ip(n1032), .op(n1053) );
  inv_1 U1489 ( .ip(n1033), .op(n1038) );
  nand2_2 U1490 ( .ip1(n1038), .ip2(n663), .op(n1044) );
  nand2_2 U1491 ( .ip1(n1042), .ip2(n1041), .op(n1043) );
  nand2_4 U1492 ( .ip1(n1044), .ip2(n1043), .op(n1438) );
  nand2_1 U1493 ( .ip1(n1438), .ip2(n1045), .op(n1051) );
  nand2_1 U1494 ( .ip1(n1890), .ip2(n1469), .op(n1049) );
  nand2_1 U1495 ( .ip1(n1896), .ip2(n1470), .op(n1048) );
  nand2_1 U1496 ( .ip1(n1888), .ip2(n1511), .op(n1047) );
  nand2_1 U1497 ( .ip1(n1893), .ip2(n1468), .op(n1046) );
  nand4_1 U1498 ( .ip1(n1049), .ip2(n1048), .ip3(n1047), .ip4(n1046), .op(
        n1422) );
  nand2_1 U1499 ( .ip1(n664), .ip2(n1506), .op(n1050) );
  nand2_1 U1500 ( .ip1(n1051), .ip2(n1050), .op(n1052) );
  nor2_1 U1501 ( .ip1(n1053), .ip2(n1052), .op(n1054) );
  nand2_1 U1502 ( .ip1(n1055), .ip2(n1054), .op(n499) );
  nand2_1 U1503 ( .ip1(n1760), .ip2(\mult/productQ [3]), .op(n1065) );
  buf_4 U1504 ( .ip(n1774), .op(n1783) );
  or2_1 U1505 ( .ip1(n1057), .ip2(n1056), .op(n1061) );
  inv_1 U1506 ( .ip(n1363), .op(n1058) );
  nand2_1 U1507 ( .ip1(n1364), .ip2(n1058), .op(n1059) );
  and2_1 U1508 ( .ip1(n1059), .ip2(n1361), .op(n1060) );
  nand2_1 U1509 ( .ip1(n1783), .ip2(n1063), .op(n1064) );
  nand2_1 U1510 ( .ip1(n1065), .ip2(n1064), .op(n486) );
  nand2_1 U1511 ( .ip1(n1067), .ip2(n1066), .op(n1068) );
  nand2_1 U1512 ( .ip1(n1760), .ip2(\mult/productQ [1]), .op(n1069) );
  nor2_1 U1513 ( .ip1(\mult/productQ [0]), .ip2(\mult/storeQ [0]), .op(n1072)
         );
  nor2_1 U1514 ( .ip1(n1072), .ip2(n1071), .op(n1073) );
  nand2_1 U1515 ( .ip1(n1783), .ip2(n1073), .op(n1075) );
  nand2_1 U1516 ( .ip1(n1760), .ip2(\mult/productQ [0]), .op(n1074) );
  inv_1 U1517 ( .ip(n1113), .op(n1077) );
  nand2_1 U1518 ( .ip1(n1802), .ip2(n1077), .op(n1079) );
  nand3_1 U1519 ( .ip1(n1078), .ip2(n1108), .ip3(n1079), .op(n1081) );
  or2_1 U1520 ( .ip1(n1079), .ip2(n1078), .op(n1080) );
  nand3_1 U1521 ( .ip1(n1082), .ip2(n1081), .ip3(n1080), .op(n1083) );
  nand2_1 U1522 ( .ip1(n573), .ip2(n1083), .op(n1085) );
  nand2_1 U1523 ( .ip1(n1085), .ip2(n1084), .op(n469) );
  nand2_1 U1524 ( .ip1(n1760), .ip2(\mult/productQ [23]), .op(n1107) );
  nor2_1 U1525 ( .ip1(n1089), .ip2(n1087), .op(n1093) );
  inv_1 U1526 ( .ip(n1089), .op(n1090) );
  nor2_1 U1527 ( .ip1(n1097), .ip2(n1108), .op(n1092) );
  nor3_2 U1528 ( .ip1(n1094), .ip2(n1093), .ip3(n1092), .op(n1099) );
  nor2_1 U1529 ( .ip1(\mult/storeQ [23]), .ip2(\mult/productQ [23]), .op(n1096) );
  and2_1 U1530 ( .ip1(\mult/productQ [23]), .ip2(\mult/storeQ [23]), .op(n1095) );
  nor2_1 U1531 ( .ip1(n1113), .ip2(n1097), .op(n1098) );
  nand2_1 U1532 ( .ip1(n1802), .ip2(n1098), .op(n1101) );
  nand3_1 U1533 ( .ip1(n1100), .ip2(n1099), .ip3(n1101), .op(n1103) );
  or2_1 U1534 ( .ip1(n1101), .ip2(n1100), .op(n1102) );
  nand3_1 U1535 ( .ip1(n1104), .ip2(n1103), .ip3(n1102), .op(n1105) );
  nand2_1 U1536 ( .ip1(n573), .ip2(n1105), .op(n1106) );
  nand2_1 U1537 ( .ip1(n1107), .ip2(n1106), .op(n466) );
  nand2_1 U1538 ( .ip1(n1760), .ip2(\mult/productQ [21]), .op(n1124) );
  nor2_1 U1539 ( .ip1(n1114), .ip2(n1108), .op(n1109) );
  nor2_1 U1540 ( .ip1(n1110), .ip2(n1109), .op(n1116) );
  nor2_1 U1541 ( .ip1(n1114), .ip2(n1113), .op(n1115) );
  nand2_1 U1542 ( .ip1(n1802), .ip2(n1115), .op(n1118) );
  nand3_1 U1543 ( .ip1(n1117), .ip2(n1116), .ip3(n1118), .op(n1120) );
  or2_1 U1544 ( .ip1(n1118), .ip2(n1117), .op(n1119) );
  nand3_1 U1545 ( .ip1(n1121), .ip2(n1120), .ip3(n1119), .op(n1122) );
  nand2_1 U1546 ( .ip1(n573), .ip2(n1122), .op(n1123) );
  nand2_1 U1547 ( .ip1(n1124), .ip2(n1123), .op(n468) );
  inv_4 U1548 ( .ip(n1852), .op(n1945) );
  nand2_1 U1549 ( .ip1(n1125), .ip2(n863), .op(n1126) );
  nand2_2 U1550 ( .ip1(n1127), .ip2(n1559), .op(n1611) );
  nor2_2 U1551 ( .ip1(n1128), .ip2(n569), .op(n1129) );
  nand2_2 U1552 ( .ip1(n1129), .ip2(n1548), .op(n1613) );
  nor2_1 U1553 ( .ip1(n1613), .ip2(n1611), .op(n1130) );
  nand2_4 U1554 ( .ip1(n1138), .ip2(result2[14]), .op(n1132) );
  nand2_4 U1555 ( .ip1(n1133), .ip2(n1132), .op(n1619) );
  nor2_2 U1556 ( .ip1(n1133), .ip2(n1132), .op(n1621) );
  nor2_2 U1557 ( .ip1(n1134), .ip2(n1621), .op(n1148) );
  nand2_1 U1558 ( .ip1(n1148), .ip2(n1135), .op(n1146) );
  nand2_1 U1559 ( .ip1(n1138), .ip2(n668), .op(n1140) );
  nand2_1 U1560 ( .ip1(n1141), .ip2(n1142), .op(n1143) );
  nand2_1 U1561 ( .ip1(n1149), .ip2(n1147), .op(n1158) );
  nor2_2 U1562 ( .ip1(n1635), .ip2(n1148), .op(n1151) );
  nand2_1 U1563 ( .ip1(n1152), .ip2(n1151), .op(n1154) );
  nand2_1 U1564 ( .ip1(n1154), .ip2(n1153), .op(n1155) );
  inv_1 U1565 ( .ip(n1155), .op(n1156) );
  nand3_1 U1566 ( .ip1(n1158), .ip2(n1157), .ip3(n1156), .op(n443) );
  nand2_1 U1567 ( .ip1(n1160), .ip2(n568), .op(n1161) );
  nand2_1 U1568 ( .ip1(n1162), .ip2(n568), .op(n1163) );
  inv_1 U1569 ( .ip(n1819), .op(n1164) );
  xor2_1 U1570 ( .ip1(n1820), .ip2(n1165), .op(n1166) );
  nand2_4 U1571 ( .ip1(n1166), .ip2(n1833), .op(n1168) );
  nand2_1 U1572 ( .ip1(n1825), .ip2(partialQ[2]), .op(n1167) );
  nor2_1 U1573 ( .ip1(n863), .ip2(n1169), .op(n1171) );
  inv_1 U1574 ( .ip(\mult/state [1]), .op(n1172) );
  nor2_2 U1575 ( .ip1(\mult/state [0]), .ip2(n1172), .op(n1849) );
  inv_1 U1576 ( .ip(n1174), .op(n1200) );
  nor2_1 U1577 ( .ip1(n1175), .ip2(n1443), .op(n1176) );
  nand2_1 U1578 ( .ip1(n966), .ip2(n1176), .op(n1187) );
  inv_1 U1579 ( .ip(n1187), .op(n1239) );
  nor2_1 U1580 ( .ip1(n1854), .ip2(n1177), .op(n1178) );
  nand2_1 U1581 ( .ip1(n1192), .ip2(n1443), .op(n1179) );
  nand2_1 U1582 ( .ip1(n1255), .ip2(n1179), .op(n1180) );
  and2_1 U1583 ( .ip1(counterD[3]), .ip2(n1181), .op(N270) );
  and2_1 U1584 ( .ip1(counterD[0]), .ip2(n1181), .op(N267) );
  and2_1 U1585 ( .ip1(counterD[1]), .ip2(n1181), .op(N268) );
  and2_1 U1586 ( .ip1(counterD[2]), .ip2(n1181), .op(N269) );
  buf_1 U1587 ( .ip(counter2Q[2]), .op(n1232) );
  nand2_1 U1588 ( .ip1(n616), .ip2(n1232), .op(n1182) );
  inv_1 U1589 ( .ip(counter2Q[0]), .op(n1225) );
  buf_1 U1590 ( .ip(counter2Q[1]), .op(n1226) );
  nand2_1 U1591 ( .ip1(n571), .ip2(n1226), .op(n1229) );
  inv_1 U1592 ( .ip(counter2Q[4]), .op(n1667) );
  and2_1 U1593 ( .ip1(n1832), .ip2(n648), .op(N287) );
  buf_1 U1594 ( .ip(counter2Q[5]), .op(n1666) );
  nand2_1 U1595 ( .ip1(n630), .ip2(n1666), .op(n1649) );
  nand2_1 U1596 ( .ip1(n578), .ip2(n617), .op(n1183) );
  nor2_1 U1597 ( .ip1(n1649), .ip2(n1183), .op(n1185) );
  inv_1 U1598 ( .ip(counter2Q[8]), .op(n1655) );
  xor2_2 U1599 ( .ip1(n1681), .ip2(n1655), .op(n1186) );
  and2_1 U1600 ( .ip1(n1832), .ip2(n1186), .op(N291) );
  nor2_2 U1601 ( .ip1(n1859), .ip2(n1858), .op(n1862) );
  nor2_1 U1602 ( .ip1(n1512), .ip2(n1187), .op(n1190) );
  nand2_1 U1603 ( .ip1(n1511), .ip2(\mult/counterQ [3]), .op(n1188) );
  nand2_1 U1604 ( .ip1(n966), .ip2(n1188), .op(n1189) );
  nand2_1 U1605 ( .ip1(n1255), .ip2(n1189), .op(n1237) );
  inv_1 U1606 ( .ip(n1191), .op(n1194) );
  nand2_1 U1607 ( .ip1(n1192), .ip2(\mult/state [1]), .op(n1193) );
  nand2_1 U1608 ( .ip1(n1194), .ip2(n1193), .op(n530) );
  inv_1 U1609 ( .ip(\mult/state [0]), .op(n1196) );
  nor3_1 U1610 ( .ip1(\mult/state [1]), .ip2(n1196), .ip3(n1195), .op(n1197)
         );
  nor3_1 U1611 ( .ip1(reset), .ip2(n1849), .ip3(n1197), .op(n528) );
  nand2_1 U1612 ( .ip1(n887), .ip2(n1198), .op(n1199) );
  nand2_1 U1613 ( .ip1(n966), .ip2(n1199), .op(n1202) );
  nand2_1 U1614 ( .ip1(n1200), .ip2(n1851), .op(n1201) );
  nand2_1 U1615 ( .ip1(n1202), .ip2(n1201), .op(n523) );
  inv_1 U1616 ( .ip(counter2Q[6]), .op(n1204) );
  nor2_1 U1617 ( .ip1(n1668), .ip2(n1649), .op(n1203) );
  and2_1 U1618 ( .ip1(n1205), .ip2(n1832), .op(N289) );
  buf_1 U1619 ( .ip(counter2Q[10]), .op(n1214) );
  inv_1 U1620 ( .ip(n1214), .op(n1207) );
  nand2_1 U1621 ( .ip1(n629), .ip2(n584), .op(n1216) );
  nor2_1 U1622 ( .ip1(n1681), .ip2(n1216), .op(n1206) );
  and2_1 U1623 ( .ip1(n1208), .ip2(n1832), .op(N293) );
  inv_1 U1624 ( .ip(n579), .op(n1212) );
  inv_1 U1625 ( .ip(n1216), .op(n1209) );
  nand2_1 U1626 ( .ip1(n1209), .ip2(n1214), .op(n1210) );
  nor2_1 U1627 ( .ip1(n1681), .ip2(n1210), .op(n1211) );
  and2_1 U1628 ( .ip1(n1213), .ip2(n1832), .op(N294) );
  inv_1 U1629 ( .ip(counter2Q[12]), .op(n1220) );
  nand2_1 U1630 ( .ip1(n579), .ip2(n1214), .op(n1215) );
  inv_1 U1631 ( .ip(n1680), .op(n1217) );
  nor2_1 U1632 ( .ip1(n1681), .ip2(n1217), .op(n1218) );
  and2_1 U1633 ( .ip1(n1219), .ip2(n1832), .op(N295) );
  inv_1 U1634 ( .ip(counter2Q[13]), .op(n1223) );
  inv_1 U1635 ( .ip(n1220), .op(n1672) );
  nand2_1 U1636 ( .ip1(n1680), .ip2(n1672), .op(n1221) );
  nor2_1 U1637 ( .ip1(n1221), .ip2(n1681), .op(n1222) );
  and2_1 U1638 ( .ip1(n1224), .ip2(n1832), .op(N296) );
  inv_1 U1639 ( .ip(n1226), .op(n1227) );
  and2_1 U1640 ( .ip1(n1832), .ip2(n1228), .op(N284) );
  inv_1 U1641 ( .ip(n1232), .op(n1230) );
  inv_1 U1642 ( .ip(n1229), .op(n1233) );
  and2_1 U1643 ( .ip1(n1832), .ip2(n1231), .op(N285) );
  and2_1 U1644 ( .ip1(n1233), .ip2(n1232), .op(n1234) );
  and2_1 U1645 ( .ip1(n1832), .ip2(n1236), .op(N286) );
  nand2_1 U1646 ( .ip1(n1237), .ip2(\mult/counterQ [5]), .op(n1241) );
  and2_1 U1647 ( .ip1(\mult/counterQ [3]), .ip2(n671), .op(n1238) );
  nand2_1 U1648 ( .ip1(n1239), .ip2(n1238), .op(n1240) );
  nand2_1 U1649 ( .ip1(n1241), .ip2(n1240), .op(n527) );
  nand2_1 U1650 ( .ip1(n1586), .ip2(state[0]), .op(n1242) );
  nor2_1 U1651 ( .ip1(n1242), .ip2(n838), .op(n1243) );
  inv_1 U1652 ( .ip(counterQ[1]), .op(n1253) );
  inv_1 U1653 ( .ip(n1253), .op(n1244) );
  inv_1 U1654 ( .ip(counterQ[2]), .op(n1251) );
  inv_1 U1655 ( .ip(n1251), .op(n1246) );
  and2_1 U1656 ( .ip1(n1245), .ip2(n1246), .op(n1247) );
  and2_1 U1657 ( .ip1(n1243), .ip2(n1249), .op(N235) );
  inv_1 U1658 ( .ip(counterQ[0]), .op(n1250) );
  and2_1 U1659 ( .ip1(n1243), .ip2(n1250), .op(N232) );
  and2_1 U1660 ( .ip1(n1243), .ip2(n1252), .op(N234) );
  and2_1 U1661 ( .ip1(n1243), .ip2(n1254), .op(N233) );
  inv_1 U1662 ( .ip(n1255), .op(n1256) );
  nand2_1 U1663 ( .ip1(n1256), .ip2(\mult/counterQ [2]), .op(n1260) );
  nand2_1 U1664 ( .ip1(n1468), .ip2(n1853), .op(n1257) );
  nand2_1 U1665 ( .ip1(n1257), .ip2(n1343), .op(n1258) );
  nand2_1 U1666 ( .ip1(n966), .ip2(n1258), .op(n1259) );
  nand2_1 U1667 ( .ip1(n1260), .ip2(n1259), .op(n524) );
  nor2_1 U1668 ( .ip1(n1264), .ip2(n1593), .op(n1267) );
  not_ab_or_c_or_d U1669 ( .ip1(n1265), .ip2(n1264), .ip3(n1635), .ip4(n1787), 
        .op(n1266) );
  or2_1 U1670 ( .ip1(n1267), .ip2(n1266), .op(n457) );
  inv_1 U1671 ( .ip(n1942), .op(n1541) );
  nor2_1 U1672 ( .ip1(n1541), .ip2(n1945), .op(n1935) );
  nor2_1 U1673 ( .ip1(n1270), .ip2(n1945), .op(n1943) );
  inv_1 U1674 ( .ip(n1907), .op(n1543) );
  nor2_1 U1675 ( .ip1(n1543), .ip2(n1945), .op(n1913) );
  nor2_1 U1676 ( .ip1(n1268), .ip2(n1945), .op(n1906) );
  nor2_1 U1677 ( .ip1(n1902), .ip2(n1268), .op(n1269) );
  nand2_1 U1678 ( .ip1(n623), .ip2(n1269), .op(n1953) );
  nor2_1 U1679 ( .ip1(n1954), .ip2(n1953), .op(n1956) );
  nand2_1 U1680 ( .ip1(n622), .ip2(n1914), .op(n1920) );
  nor2_1 U1681 ( .ip1(n1917), .ip2(n1920), .op(n1919) );
  nor2_1 U1682 ( .ip1(n1944), .ip2(n1270), .op(n1271) );
  nand2_1 U1683 ( .ip1(n623), .ip2(n1271), .op(n1949) );
  nor2_1 U1684 ( .ip1(n1950), .ip2(n1949), .op(n1952) );
  nand2_1 U1685 ( .ip1(n622), .ip2(n1926), .op(n1929) );
  nor2_1 U1686 ( .ip1(n1930), .ip2(n1929), .op(n1932) );
  inv_1 U1687 ( .ip(n1272), .op(n1273) );
  nand2_1 U1688 ( .ip1(n1825), .ip2(partialQ[4]), .op(n1275) );
  nand2_1 U1689 ( .ip1(n1276), .ip2(n1275), .op(n453) );
  nor2_1 U1690 ( .ip1(n1319), .ip2(n1342), .op(n1278) );
  nor2_1 U1691 ( .ip1(n1317), .ip2(n1406), .op(n1277) );
  nor2_1 U1692 ( .ip1(n1278), .ip2(n1277), .op(n1282) );
  nor2_1 U1693 ( .ip1(n1343), .ip2(n1318), .op(n1280) );
  nor2_1 U1694 ( .ip1(n1443), .ip2(n1316), .op(n1279) );
  nor2_1 U1695 ( .ip1(n1280), .ip2(n1279), .op(n1281) );
  nand2_1 U1696 ( .ip1(n1282), .ip2(n1281), .op(n1418) );
  nand2_1 U1697 ( .ip1(n1519), .ip2(\mult/storeQ [23]), .op(n1289) );
  nand2_1 U1698 ( .ip1(n1889), .ip2(n1511), .op(n1287) );
  nand2_1 U1699 ( .ip1(n1891), .ip2(n1469), .op(n1286) );
  nand2_1 U1700 ( .ip1(n1894), .ip2(n1468), .op(n1285) );
  nand2_1 U1701 ( .ip1(n1897), .ip2(n1470), .op(n1284) );
  nand4_1 U1702 ( .ip1(n1287), .ip2(n1286), .ip3(n1285), .ip4(n1284), .op(
        n1417) );
  nand2_1 U1703 ( .ip1(n655), .ip2(n1417), .op(n1288) );
  nand3_1 U1704 ( .ip1(n1290), .ip2(n1289), .ip3(n1288), .op(n498) );
  nand2_1 U1705 ( .ip1(n1548), .ip2(n635), .op(n1299) );
  nor2_1 U1706 ( .ip1(n1635), .ip2(n1299), .op(n1298) );
  nand2_1 U1707 ( .ip1(n631), .ip2(n659), .op(n1305) );
  nand2_1 U1708 ( .ip1(n631), .ip2(n603), .op(n1300) );
  nand4_1 U1709 ( .ip1(n1301), .ip2(n1298), .ip3(n1305), .ip4(n1300), .op(
        n1311) );
  nand2_1 U1710 ( .ip1(n1299), .ip2(n1833), .op(n1306) );
  nor2_1 U1711 ( .ip1(n1306), .ip2(n1300), .op(n1303) );
  nor2_1 U1712 ( .ip1(n1306), .ip2(n1301), .op(n1302) );
  nor2_1 U1713 ( .ip1(n1303), .ip2(n1302), .op(n1310) );
  nor2_1 U1714 ( .ip1(n1304), .ip2(n1593), .op(n1308) );
  nor2_1 U1715 ( .ip1(n1306), .ip2(n1305), .op(n1307) );
  nor2_1 U1716 ( .ip1(n1308), .ip2(n1307), .op(n1309) );
  nand3_1 U1717 ( .ip1(n1309), .ip2(n1310), .ip3(n1311), .op(n449) );
  nor2_1 U1718 ( .ip1(n1317), .ip2(n1318), .op(n1313) );
  nor2_1 U1719 ( .ip1(n1319), .ip2(n1316), .op(n1312) );
  inv_1 U1720 ( .ip(n1347), .op(n1402) );
  nand2_1 U1721 ( .ip1(n1438), .ip2(n1402), .op(n1315) );
  nand2_1 U1722 ( .ip1(n1519), .ip2(\mult/storeQ [3]), .op(n1314) );
  nand2_1 U1723 ( .ip1(n1315), .ip2(n1314), .op(n518) );
  nor2_1 U1724 ( .ip1(n1343), .ip2(n1316), .op(n1322) );
  nor2_1 U1725 ( .ip1(n1317), .ip2(n1342), .op(n1321) );
  nor2_1 U1726 ( .ip1(n1319), .ip2(n1318), .op(n1320) );
  nor3_2 U1727 ( .ip1(n1322), .ip2(n1321), .ip3(n1320), .op(n1507) );
  inv_1 U1728 ( .ip(n1507), .op(n1413) );
  nand2_1 U1729 ( .ip1(n1438), .ip2(n1413), .op(n1324) );
  nand2_1 U1730 ( .ip1(n1519), .ip2(\mult/storeQ [5]), .op(n1323) );
  nand2_1 U1731 ( .ip1(n1324), .ip2(n1323), .op(n516) );
  nor2_1 U1732 ( .ip1(n1874), .ip2(\mult/counterQ [2]), .op(n1325) );
  nand2_1 U1733 ( .ip1(n1880), .ip2(n1325), .op(n1326) );
  inv_1 U1734 ( .ip(n1326), .op(n1476) );
  nand2_1 U1735 ( .ip1(n1438), .ip2(n1476), .op(n1328) );
  nand2_1 U1736 ( .ip1(n1519), .ip2(\mult/storeQ [0]), .op(n1327) );
  nand2_1 U1737 ( .ip1(n1328), .ip2(n1327), .op(n521) );
  nand2_1 U1738 ( .ip1(n1882), .ip2(n1892), .op(n1330) );
  nand2_1 U1739 ( .ip1(n1883), .ip2(n1470), .op(n1329) );
  nand2_1 U1740 ( .ip1(n1438), .ip2(n1461), .op(n1332) );
  nand2_1 U1741 ( .ip1(n1519), .ip2(\mult/storeQ [2]), .op(n1331) );
  nand2_1 U1742 ( .ip1(n1332), .ip2(n1331), .op(n519) );
  nand2_1 U1743 ( .ip1(n1883), .ip2(n1468), .op(n1334) );
  nand2_1 U1744 ( .ip1(n1886), .ip2(n1470), .op(n1333) );
  nand2_1 U1745 ( .ip1(n1438), .ip2(n1449), .op(n1336) );
  nand2_1 U1746 ( .ip1(n1519), .ip2(\mult/storeQ [4]), .op(n1335) );
  nand2_1 U1747 ( .ip1(n1336), .ip2(n1335), .op(n517) );
  nand2_1 U1748 ( .ip1(n1438), .ip2(n1386), .op(n1338) );
  nand2_1 U1749 ( .ip1(n1480), .ip2(\mult/storeQ [1]), .op(n1337) );
  nand2_1 U1750 ( .ip1(n1338), .ip2(n1337), .op(n520) );
  nand2_1 U1751 ( .ip1(n1889), .ip2(n1468), .op(n1340) );
  nand2_1 U1752 ( .ip1(n1891), .ip2(n1470), .op(n1339) );
  nor2_1 U1753 ( .ip1(n1443), .ip2(n1342), .op(n1345) );
  nor2_1 U1754 ( .ip1(n1343), .ip2(n1406), .op(n1344) );
  nor2_1 U1755 ( .ip1(n1345), .ip2(n1344), .op(n1346) );
  nand2_1 U1756 ( .ip1(n1341), .ip2(n1346), .op(n1401) );
  nor2_1 U1757 ( .ip1(n1034), .ip2(n1347), .op(n1348) );
  nand2_1 U1758 ( .ip1(n1283), .ip2(n1348), .op(n1355) );
  mux2_4 U1759 ( .ip1(n1897), .ip2(n1894), .s(n1349), .op(n1350) );
  nand2_1 U1760 ( .ip1(n1350), .ip2(\mult/counterQ [2]), .op(n1351) );
  nor2_1 U1761 ( .ip1(\mult/counterQ [3]), .ip2(n1351), .op(n1352) );
  nand2_1 U1762 ( .ip1(n607), .ip2(n1352), .op(n1354) );
  nand4_1 U1763 ( .ip1(n1356), .ip2(n1355), .ip3(n1354), .ip4(n1353), .op(n502) );
  nand2_1 U1764 ( .ip1(n1760), .ip2(\mult/productQ [4]), .op(n1360) );
  nand2_1 U1765 ( .ip1(n1696), .ip2(n1698), .op(n1357) );
  xnor2_2 U1766 ( .ip1(n1357), .ip2(n1697), .op(n1358) );
  nand2_1 U1767 ( .ip1(n1783), .ip2(n1358), .op(n1359) );
  nand2_1 U1768 ( .ip1(n1360), .ip2(n1359), .op(n485) );
  nand2_1 U1769 ( .ip1(n1760), .ip2(\mult/productQ [2]), .op(n1368) );
  inv_1 U1770 ( .ip(n1361), .op(n1362) );
  or2_1 U1771 ( .ip1(n1363), .ip2(n1362), .op(n1365) );
  xnor2_2 U1772 ( .ip1(n1365), .ip2(n1364), .op(n1366) );
  nand2_1 U1773 ( .ip1(n1783), .ip2(n1366), .op(n1367) );
  nand2_1 U1774 ( .ip1(n1368), .ip2(n1367), .op(n487) );
  nand2_1 U1775 ( .ip1(n1760), .ip2(\mult/productQ [7]), .op(n1383) );
  nand2_1 U1776 ( .ip1(n1371), .ip2(n1374), .op(n1373) );
  inv_1 U1777 ( .ip(n1778), .op(n1372) );
  inv_1 U1778 ( .ip(n1375), .op(n1376) );
  nand2_1 U1779 ( .ip1(n1697), .ip2(n1376), .op(n1780) );
  nor2_1 U1780 ( .ip1(n1777), .ip2(n1780), .op(n1377) );
  nor2_1 U1781 ( .ip1(n1378), .ip2(n1377), .op(n1379) );
  xor2_1 U1782 ( .ip1(n1380), .ip2(n1379), .op(n1381) );
  nand2_4 U1783 ( .ip1(n1381), .ip2(n1810), .op(n1382) );
  nand2_1 U1784 ( .ip1(n1383), .ip2(n1382), .op(n482) );
  inv_1 U1785 ( .ip(n1384), .op(n1385) );
  nand2_1 U1786 ( .ip1(n1387), .ip2(n607), .op(n1389) );
  nand2_1 U1787 ( .ip1(n1480), .ip2(\mult/storeQ [9]), .op(n1388) );
  nand2_1 U1788 ( .ip1(n1389), .ip2(n1388), .op(n512) );
  nand2_1 U1789 ( .ip1(n1438), .ip2(n1418), .op(n1391) );
  nand2_1 U1790 ( .ip1(n1480), .ip2(\mult/storeQ [7]), .op(n1390) );
  nand2_1 U1791 ( .ip1(n1391), .ip2(n1390), .op(n514) );
  nand2_1 U1792 ( .ip1(n1438), .ip2(n1423), .op(n1393) );
  nand2_1 U1793 ( .ip1(n1480), .ip2(\mult/storeQ [6]), .op(n1392) );
  nand2_1 U1794 ( .ip1(n1393), .ip2(n1392), .op(n515) );
  nand2_1 U1795 ( .ip1(n1887), .ip2(n1468), .op(n1397) );
  nand2_1 U1796 ( .ip1(n1888), .ip2(n1470), .op(n1396) );
  nand2_1 U1797 ( .ip1(n1883), .ip2(n1511), .op(n1395) );
  nand2_1 U1798 ( .ip1(n1886), .ip2(n1469), .op(n1394) );
  nand2_1 U1799 ( .ip1(n1438), .ip2(n1467), .op(n1400) );
  nand2_1 U1800 ( .ip1(n655), .ip2(n1476), .op(n1399) );
  nand2_1 U1801 ( .ip1(n1519), .ip2(\mult/storeQ [8]), .op(n1398) );
  nand3_1 U1802 ( .ip1(n1400), .ip2(n1399), .ip3(n1398), .op(n513) );
  nand2_1 U1803 ( .ip1(n1438), .ip2(n1401), .op(n1405) );
  nand2_1 U1804 ( .ip1(n655), .ip2(n1402), .op(n1404) );
  nand2_1 U1805 ( .ip1(n1480), .ip2(\mult/storeQ [11]), .op(n1403) );
  nand3_1 U1806 ( .ip1(n1405), .ip2(n1404), .ip3(n1403), .op(n510) );
  and2_1 U1807 ( .ip1(n1894), .ip2(n955), .op(n1411) );
  nor2_1 U1808 ( .ip1(n1443), .ip2(n1406), .op(n1410) );
  nand2_1 U1809 ( .ip1(n1889), .ip2(n1469), .op(n1408) );
  nand2_1 U1810 ( .ip1(n1891), .ip2(n1468), .op(n1407) );
  nand2_1 U1811 ( .ip1(n1408), .ip2(n1407), .op(n1409) );
  nor3_2 U1812 ( .ip1(n1411), .ip2(n1410), .ip3(n1409), .op(n1509) );
  inv_1 U1813 ( .ip(n1509), .op(n1412) );
  nand2_1 U1814 ( .ip1(n1438), .ip2(n1412), .op(n1416) );
  nand2_1 U1815 ( .ip1(n655), .ip2(n1413), .op(n1415) );
  nand2_1 U1816 ( .ip1(n1480), .ip2(\mult/storeQ [13]), .op(n1414) );
  nand3_1 U1817 ( .ip1(n1416), .ip2(n1415), .ip3(n1414), .op(n508) );
  nand2_1 U1818 ( .ip1(n1438), .ip2(n1417), .op(n1421) );
  nand2_1 U1819 ( .ip1(n655), .ip2(n1418), .op(n1420) );
  nand2_1 U1820 ( .ip1(n1480), .ip2(\mult/storeQ [15]), .op(n1419) );
  nand3_1 U1821 ( .ip1(n1421), .ip2(n1420), .ip3(n1419), .op(n506) );
  nand2_1 U1822 ( .ip1(n1438), .ip2(n1422), .op(n1426) );
  nand2_1 U1823 ( .ip1(n655), .ip2(n1423), .op(n1425) );
  nand2_1 U1824 ( .ip1(n1480), .ip2(\mult/storeQ [14]), .op(n1424) );
  nand3_1 U1825 ( .ip1(n1426), .ip2(n1425), .ip3(n1424), .op(n507) );
  nand2_1 U1826 ( .ip1(n1888), .ip2(n1469), .op(n1430) );
  nand2_1 U1827 ( .ip1(n1893), .ip2(n1470), .op(n1429) );
  nand2_1 U1828 ( .ip1(n1887), .ip2(n1511), .op(n1428) );
  nand2_1 U1829 ( .ip1(n1890), .ip2(n1468), .op(n1427) );
  nand2_1 U1830 ( .ip1(n1438), .ip2(n1442), .op(n1433) );
  nand2_1 U1831 ( .ip1(n655), .ip2(n1449), .op(n1432) );
  nand2_1 U1832 ( .ip1(n1480), .ip2(\mult/storeQ [12]), .op(n1431) );
  nand3_1 U1833 ( .ip1(n1433), .ip2(n1432), .ip3(n1431), .op(n509) );
  nand2_1 U1834 ( .ip1(n1888), .ip2(n1468), .op(n1437) );
  nand2_1 U1835 ( .ip1(n1890), .ip2(n1470), .op(n1436) );
  nand2_1 U1836 ( .ip1(n1886), .ip2(n1511), .op(n1435) );
  nand2_1 U1837 ( .ip1(n1887), .ip2(n1469), .op(n1434) );
  nand2_1 U1838 ( .ip1(n1438), .ip2(n1455), .op(n1441) );
  nand2_1 U1839 ( .ip1(n655), .ip2(n1461), .op(n1440) );
  nand2_1 U1840 ( .ip1(n1480), .ip2(\mult/storeQ [10]), .op(n1439) );
  nand3_1 U1841 ( .ip1(n1441), .ip2(n1440), .ip3(n1439), .op(n511) );
  inv_1 U1842 ( .ip(n1442), .op(n1451) );
  nand2_1 U1843 ( .ip1(n1895), .ip2(\mult/counterQ [2]), .op(n1444) );
  and2_1 U1844 ( .ip1(n1444), .ip2(n1443), .op(n1447) );
  nor2_1 U1845 ( .ip1(n1445), .ip2(n1896), .op(n1446) );
  nand2_1 U1846 ( .ip1(n1452), .ip2(n1518), .op(n1454) );
  nand2_1 U1847 ( .ip1(n1519), .ip2(\mult/storeQ [20]), .op(n1453) );
  nand2_1 U1848 ( .ip1(n1453), .ip2(n1454), .op(n501) );
  inv_1 U1849 ( .ip(n1455), .op(n1463) );
  nand2_1 U1850 ( .ip1(n1456), .ip2(n1892), .op(n1459) );
  nand2_1 U1851 ( .ip1(n1893), .ip2(n1511), .op(n1458) );
  nand2_1 U1852 ( .ip1(n1896), .ip2(n1469), .op(n1457) );
  nor2_1 U1853 ( .ip1(n1461), .ip2(n1506), .op(n1462) );
  nand2_1 U1854 ( .ip1(n1480), .ip2(\mult/storeQ [18]), .op(n1465) );
  nand2_1 U1855 ( .ip1(n1466), .ip2(n1465), .op(n503) );
  inv_1 U1856 ( .ip(n1467), .op(n1478) );
  nand2_1 U1857 ( .ip1(n1896), .ip2(n1468), .op(n1474) );
  nand2_1 U1858 ( .ip1(n1893), .ip2(n1469), .op(n1473) );
  nand2_1 U1859 ( .ip1(n1890), .ip2(n1511), .op(n1472) );
  nand2_1 U1860 ( .ip1(n1895), .ip2(n1470), .op(n1471) );
  nor2_1 U1861 ( .ip1(n1476), .ip2(n1506), .op(n1477) );
  nand2_1 U1862 ( .ip1(n1480), .ip2(\mult/storeQ [16]), .op(n1481) );
  nand2_1 U1863 ( .ip1(n1482), .ip2(n1481), .op(n505) );
  nor2_2 U1864 ( .ip1(n1635), .ip2(n1493), .op(n1488) );
  nand2_1 U1865 ( .ip1(n1485), .ip2(n1488), .op(n1498) );
  nor2_1 U1866 ( .ip1(n1486), .ip2(n1593), .op(n1491) );
  inv_1 U1867 ( .ip(n1488), .op(n1489) );
  nor2_1 U1868 ( .ip1(n1492), .ip2(n1489), .op(n1490) );
  nor2_1 U1869 ( .ip1(n1491), .ip2(n1490), .op(n1497) );
  and3_1 U1870 ( .ip1(n1493), .ip2(n1492), .ip3(n1833), .op(n1494) );
  nand2_1 U1871 ( .ip1(n1495), .ip2(n1494), .op(n1496) );
  nand3_1 U1872 ( .ip1(n1498), .ip2(n1497), .ip3(n1496), .op(n451) );
  nand2_1 U1873 ( .ip1(n1767), .ip2(n1708), .op(n1500) );
  nand2_1 U1874 ( .ip1(n1500), .ip2(n1711), .op(n1501) );
  xor2_1 U1875 ( .ip1(n1502), .ip2(n1501), .op(n1503) );
  nand2_4 U1876 ( .ip1(n1503), .ip2(n1810), .op(n1505) );
  nand2_1 U1877 ( .ip1(n1760), .ip2(\mult/productQ [10]), .op(n1504) );
  nand2_1 U1878 ( .ip1(n1505), .ip2(n1504), .op(n479) );
  inv_1 U1879 ( .ip(n1506), .op(n1508) );
  nand2_1 U1880 ( .ip1(n1508), .ip2(n1507), .op(n1517) );
  nand2_1 U1881 ( .ip1(n1509), .ip2(n1034), .op(n1510) );
  nand2_1 U1882 ( .ip1(n1510), .ip2(n539), .op(n1515) );
  and2_1 U1883 ( .ip1(n1897), .ip2(n1511), .op(n1513) );
  nand2_1 U1884 ( .ip1(n1513), .ip2(n1512), .op(n1514) );
  nand2_1 U1885 ( .ip1(n1515), .ip2(n1514), .op(n1516) );
  nand2_1 U1886 ( .ip1(n1519), .ip2(\mult/storeQ [21]), .op(n1520) );
  nand2_1 U1887 ( .ip1(n1523), .ip2(n1522), .op(n1524) );
  inv_1 U1888 ( .ip(n1527), .op(n1528) );
  nor2_1 U1889 ( .ip1(n1635), .ip2(n1532), .op(n1530) );
  nand2_1 U1890 ( .ip1(n1531), .ip2(n1530), .op(n1540) );
  inv_1 U1891 ( .ip(n1532), .op(n1536) );
  nor3_1 U1892 ( .ip1(n604), .ip2(n1635), .ip3(n1536), .op(n1533) );
  nand2_1 U1893 ( .ip1(n1534), .ip2(n1533), .op(n1539) );
  nand2_1 U1894 ( .ip1(n1825), .ip2(partialQ[5]), .op(n1538) );
  nand3_1 U1895 ( .ip1(n1536), .ip2(n1833), .ip3(n604), .op(n1537) );
  nand4_1 U1896 ( .ip1(n1540), .ip2(n1539), .ip3(n1538), .ip4(n1537), .op(n452) );
  inv_1 U1897 ( .ip(n1921), .op(n6) );
  inv_1 U1898 ( .ip(n1948), .op(n15) );
  inv_1 U1899 ( .ip(n1904), .op(n1) );
  inv_1 U1900 ( .ip(n1928), .op(n10) );
  nand2_1 U1901 ( .ip1(n622), .ip2(n1541), .op(n1542) );
  nand2_1 U1902 ( .ip1(n1542), .ip2(n1544), .op(n1936) );
  nor2_1 U1903 ( .ip1(n1937), .ip2(n1936), .op(n1938) );
  inv_1 U1904 ( .ip(n1940), .op(n13) );
  nand2_1 U1905 ( .ip1(n623), .ip2(n1543), .op(n1545) );
  nand2_1 U1906 ( .ip1(n1545), .ip2(n1544), .op(n1912) );
  nor2_1 U1907 ( .ip1(n1908), .ip2(n1912), .op(n1909) );
  inv_1 U1908 ( .ip(n1911), .op(n3) );
  nand2_1 U1909 ( .ip1(n1587), .ip2(n633), .op(n1552) );
  nand2_1 U1910 ( .ip1(n614), .ip2(n660), .op(n1547) );
  nand2_1 U1911 ( .ip1(n1825), .ip2(partialQ[10]), .op(n1546) );
  nand2_1 U1912 ( .ip1(n567), .ip2(n1548), .op(n1588) );
  inv_1 U1913 ( .ip(n1588), .op(n1551) );
  and2_1 U1914 ( .ip1(n1551), .ip2(n660), .op(n1550) );
  nand2_1 U1915 ( .ip1(n626), .ip2(n1551), .op(n1554) );
  nor3_1 U1916 ( .ip1(n1635), .ip2(n614), .ip3(n1552), .op(n1553) );
  nand2_1 U1917 ( .ip1(n1554), .ip2(n1553), .op(n1555) );
  nand2_1 U1918 ( .ip1(n1556), .ip2(n1555), .op(n447) );
  inv_1 U1919 ( .ip(n1613), .op(n1557) );
  nand2_1 U1920 ( .ip1(n1614), .ip2(n1557), .op(n1562) );
  buf_1 U1921 ( .ip(n1618), .op(n1567) );
  inv_1 U1922 ( .ip(n605), .op(n1565) );
  nor2_2 U1923 ( .ip1(n1635), .ip2(n1564), .op(n1568) );
  or2_1 U1924 ( .ip1(n1566), .ip2(n1593), .op(n1570) );
  nand2_1 U1925 ( .ip1(n1567), .ip2(n1568), .op(n1569) );
  and2_1 U1926 ( .ip1(n1570), .ip2(n1569), .op(n1571) );
  inv_1 U1927 ( .ip(n1688), .op(n1576) );
  nand2_1 U1928 ( .ip1(n1802), .ip2(n1576), .op(n1577) );
  nand2_1 U1929 ( .ip1(n1577), .ip2(n1686), .op(n1578) );
  nand2_1 U1930 ( .ip1(n1760), .ip2(\mult/productQ [17]), .op(n1580) );
  nand2_1 U1931 ( .ip1(n1581), .ip2(n1580), .op(n472) );
  nand2_1 U1932 ( .ip1(n1802), .ip2(n1799), .op(n1582) );
  nand2_1 U1933 ( .ip1(n1582), .ip2(n1803), .op(n1583) );
  nand2_1 U1934 ( .ip1(n1760), .ip2(\mult/productQ [18]), .op(n1585) );
  nor2_1 U1935 ( .ip1(state[0]), .ip2(n1586), .op(n532) );
  inv_1 U1936 ( .ip(n1587), .op(n1596) );
  nor2_1 U1937 ( .ip1(n1596), .ip2(n1588), .op(n1589) );
  nor2_1 U1938 ( .ip1(n1591), .ip2(n1590), .op(n1604) );
  nor2_1 U1939 ( .ip1(n1635), .ip2(n1604), .op(n1595) );
  nor2_1 U1940 ( .ip1(n1594), .ip2(n1593), .op(n1603) );
  inv_1 U1941 ( .ip(n1595), .op(n1601) );
  inv_1 U1942 ( .ip(n1596), .op(n1597) );
  nand2_1 U1943 ( .ip1(n1597), .ip2(n614), .op(n1598) );
  nand2_1 U1944 ( .ip1(n633), .ip2(n1598), .op(n1605) );
  inv_1 U1945 ( .ip(n1605), .op(n1600) );
  nor2_1 U1946 ( .ip1(n1603), .ip2(n1602), .op(n1609) );
  nand2_1 U1947 ( .ip1(n1604), .ip2(n1833), .op(n1606) );
  nor2_1 U1948 ( .ip1(n1606), .ip2(n1605), .op(n1607) );
  nand2_1 U1949 ( .ip1(n1607), .ip2(n606), .op(n1608) );
  nand3_1 U1950 ( .ip1(n1608), .ip2(n1609), .ip3(n1610), .op(n446) );
  inv_2 U1951 ( .ip(n1611), .op(n1612) );
  nor2_1 U1952 ( .ip1(n1613), .ip2(n1616), .op(n1615) );
  nand2_1 U1953 ( .ip1(n1639), .ip2(n1629), .op(n1630) );
  inv_1 U1954 ( .ip(n1630), .op(n1631) );
  nand2_1 U1955 ( .ip1(n1632), .ip2(n1631), .op(n1648) );
  inv_1 U1956 ( .ip(n1632), .op(n1636) );
  nor2_2 U1957 ( .ip1(n1635), .ip2(n666), .op(n1642) );
  nand2_1 U1958 ( .ip1(n1636), .ip2(n1642), .op(n1647) );
  nand2_1 U1959 ( .ip1(n1640), .ip2(n1639), .op(n1641) );
  nand2_1 U1960 ( .ip1(n1641), .ip2(n1642), .op(n1643) );
  nand2_1 U1961 ( .ip1(n1644), .ip2(n1643), .op(n1645) );
  inv_1 U1962 ( .ip(n1645), .op(n1646) );
  nand3_1 U1963 ( .ip1(n1648), .ip2(n1647), .ip3(n1646), .op(n442) );
  inv_1 U1964 ( .ip(n578), .op(n1653) );
  inv_1 U1965 ( .ip(n1649), .op(n1650) );
  nand2_1 U1966 ( .ip1(n1650), .ip2(n617), .op(n1651) );
  and2_1 U1967 ( .ip1(n1654), .ip2(n1832), .op(N290) );
  inv_1 U1968 ( .ip(counter2Q[9]), .op(n1657) );
  and2_1 U1969 ( .ip1(n1658), .ip2(n1832), .op(N292) );
  nand2_1 U1970 ( .ip1(n1760), .ip2(\mult/productQ [8]), .op(n1665) );
  inv_1 U1971 ( .ip(n1659), .op(n1660) );
  xor2_1 U1972 ( .ip1(n1662), .ip2(n1767), .op(n1663) );
  nand2_4 U1973 ( .ip1(n1663), .ip2(n1810), .op(n1664) );
  nand2_1 U1974 ( .ip1(n1665), .ip2(n1664), .op(n481) );
  inv_1 U1975 ( .ip(n1666), .op(n1670) );
  and2_1 U1976 ( .ip1(n1671), .ip2(n1832), .op(N288) );
  inv_1 U1977 ( .ip(counter2Q[15]), .op(n1676) );
  nand2_1 U1978 ( .ip1(n585), .ip2(n1672), .op(n1678) );
  inv_1 U1979 ( .ip(counter2Q[14]), .op(n1684) );
  nor2_1 U1980 ( .ip1(n1678), .ip2(n1684), .op(n1673) );
  nand2_1 U1981 ( .ip1(n1680), .ip2(n1673), .op(n1674) );
  nor2_1 U1982 ( .ip1(n1674), .ip2(n1681), .op(n1675) );
  and2_1 U1983 ( .ip1(n1677), .ip2(n1832), .op(N298) );
  inv_1 U1984 ( .ip(n1678), .op(n1679) );
  nand2_1 U1985 ( .ip1(n1680), .ip2(n1679), .op(n1682) );
  nor2_1 U1986 ( .ip1(n1682), .ip2(n1681), .op(n1683) );
  and2_1 U1987 ( .ip1(n1685), .ip2(n1832), .op(N297) );
  inv_1 U1988 ( .ip(n1686), .op(n1687) );
  nor2_1 U1989 ( .ip1(n1688), .ip2(n1687), .op(n1689) );
  xor2_1 U1990 ( .ip1(n1689), .ip2(n1802), .op(n1690) );
  nand2_4 U1991 ( .ip1(n1690), .ip2(n1783), .op(n1692) );
  nand2_1 U1992 ( .ip1(n1760), .ip2(\mult/productQ [16]), .op(n1691) );
  nand2_1 U1993 ( .ip1(n1692), .ip2(n1691), .op(n473) );
  nand2_1 U1994 ( .ip1(n1760), .ip2(\mult/productQ [5]), .op(n1704) );
  or2_1 U1995 ( .ip1(n1695), .ip2(n1694), .op(n1701) );
  nand2_1 U1996 ( .ip1(n1697), .ip2(n1696), .op(n1699) );
  nand2_1 U1997 ( .ip1(n1699), .ip2(n1698), .op(n1700) );
  xnor2_1 U1998 ( .ip1(n1701), .ip2(n1700), .op(n1702) );
  nand2_1 U1999 ( .ip1(n1704), .ip2(n1703), .op(n484) );
  inv_1 U2000 ( .ip(n1705), .op(n1706) );
  inv_1 U2001 ( .ip(n1708), .op(n1709) );
  nor2_1 U2002 ( .ip1(n1712), .ip2(n1709), .op(n1710) );
  nand2_1 U2003 ( .ip1(n1767), .ip2(n1710), .op(n1716) );
  nor2_1 U2004 ( .ip1(n1712), .ip2(n1711), .op(n1713) );
  nor2_1 U2005 ( .ip1(n1714), .ip2(n1713), .op(n1715) );
  nand2_1 U2006 ( .ip1(n1716), .ip2(n1715), .op(n1717) );
  xor2_1 U2007 ( .ip1(n1718), .ip2(n1717), .op(n1719) );
  nand2_4 U2008 ( .ip1(n1719), .ip2(n1783), .op(n1721) );
  nand2_1 U2009 ( .ip1(n1760), .ip2(\mult/productQ [11]), .op(n1720) );
  nand2_1 U2010 ( .ip1(n1721), .ip2(n1720), .op(n478) );
  inv_1 U2011 ( .ip(n1722), .op(n1723) );
  nor2_1 U2012 ( .ip1(n1724), .ip2(n1723), .op(n1730) );
  nor2_1 U2013 ( .ip1(n1764), .ip2(n1765), .op(n1725) );
  nand2_1 U2014 ( .ip1(n1767), .ip2(n1725), .op(n1728) );
  nor2_1 U2015 ( .ip1(n1764), .ip2(n1768), .op(n1726) );
  nor2_1 U2016 ( .ip1(n1763), .ip2(n1726), .op(n1727) );
  nand2_1 U2017 ( .ip1(n1728), .ip2(n1727), .op(n1729) );
  xor2_1 U2018 ( .ip1(n1730), .ip2(n1729), .op(n1731) );
  nand2_1 U2019 ( .ip1(n1760), .ip2(\mult/productQ [13]), .op(n1732) );
  inv_1 U2020 ( .ip(n1750), .op(n1733) );
  nor2_1 U2021 ( .ip1(n1745), .ip2(n1733), .op(n1740) );
  inv_1 U2022 ( .ip(n1746), .op(n1735) );
  nor2_1 U2023 ( .ip1(n1735), .ip2(n1765), .op(n1734) );
  nand2_1 U2024 ( .ip1(n1767), .ip2(n1734), .op(n1738) );
  nor2_1 U2025 ( .ip1(n1735), .ip2(n1768), .op(n1736) );
  nand2_1 U2026 ( .ip1(n1738), .ip2(n1737), .op(n1739) );
  xor2_1 U2027 ( .ip1(n1740), .ip2(n1739), .op(n1741) );
  nand2_1 U2028 ( .ip1(n1760), .ip2(\mult/productQ [14]), .op(n1742) );
  inv_1 U2029 ( .ip(n1745), .op(n1748) );
  nand2_1 U2030 ( .ip1(n1746), .ip2(n1748), .op(n1752) );
  nor2_1 U2031 ( .ip1(n1752), .ip2(n1765), .op(n1747) );
  nand2_1 U2032 ( .ip1(n1767), .ip2(n1747), .op(n1756) );
  nand2_1 U2033 ( .ip1(n1749), .ip2(n1748), .op(n1751) );
  nand2_1 U2034 ( .ip1(n1751), .ip2(n1750), .op(n1754) );
  nor2_1 U2035 ( .ip1(n1752), .ip2(n1768), .op(n1753) );
  nand2_1 U2036 ( .ip1(n1756), .ip2(n1755), .op(n1757) );
  xor2_1 U2037 ( .ip1(n1758), .ip2(n1757), .op(n1759) );
  nand2_4 U2038 ( .ip1(n1759), .ip2(n1810), .op(n1762) );
  nand2_1 U2039 ( .ip1(n1760), .ip2(\mult/productQ [15]), .op(n1761) );
  nand2_1 U2040 ( .ip1(n1762), .ip2(n1761), .op(n474) );
  nor2_1 U2041 ( .ip1(n1764), .ip2(n1763), .op(n1771) );
  inv_1 U2042 ( .ip(n1765), .op(n1766) );
  nand2_1 U2043 ( .ip1(n1767), .ip2(n1766), .op(n1769) );
  nand2_1 U2044 ( .ip1(n1769), .ip2(n1768), .op(n1770) );
  nand2_1 U2045 ( .ip1(n573), .ip2(n1773), .op(n1776) );
  nand2_1 U2046 ( .ip1(n1760), .ip2(\mult/productQ [12]), .op(n1775) );
  nand2_1 U2047 ( .ip1(n1776), .ip2(n1775), .op(n477) );
  nand2_1 U2048 ( .ip1(n1760), .ip2(\mult/productQ [6]), .op(n1786) );
  nand2_1 U2049 ( .ip1(n1780), .ip2(n1779), .op(n1781) );
  xor2_1 U2050 ( .ip1(n1782), .ip2(n1781), .op(n1784) );
  nand2_4 U2051 ( .ip1(n1784), .ip2(n1810), .op(n1785) );
  nand2_1 U2052 ( .ip1(n1786), .ip2(n1785), .op(n483) );
  nor2_1 U2053 ( .ip1(n571), .ip2(n642), .op(N283) );
  nand2_1 U2054 ( .ip1(n1789), .ip2(n647), .op(n1790) );
  nand2_1 U2055 ( .ip1(n1791), .ip2(n1790), .op(n1792) );
  xor2_1 U2056 ( .ip1(n1263), .ip2(n1792), .op(n1793) );
  nand2_4 U2057 ( .ip1(n1793), .ip2(n1833), .op(n1795) );
  nand2_1 U2058 ( .ip1(n1825), .ip2(partialQ[1]), .op(n1794) );
  nand2_1 U2059 ( .ip1(n1795), .ip2(n1794), .op(n456) );
  inv_1 U2060 ( .ip(n1796), .op(n1797) );
  inv_1 U2061 ( .ip(n1799), .op(n1800) );
  nor2_1 U2062 ( .ip1(n1804), .ip2(n1800), .op(n1801) );
  nand2_1 U2063 ( .ip1(n1802), .ip2(n1801), .op(n1808) );
  nor2_1 U2064 ( .ip1(n1804), .ip2(n1803), .op(n1805) );
  nor2_1 U2065 ( .ip1(n1806), .ip2(n1805), .op(n1807) );
  nand2_1 U2066 ( .ip1(n1808), .ip2(n1807), .op(n1809) );
  nand2_1 U2067 ( .ip1(n1760), .ip2(\mult/productQ [19]), .op(n1812) );
  nand2_1 U2068 ( .ip1(n1813), .ip2(n1812), .op(n470) );
  nand2_1 U2069 ( .ip1(n738), .ip2(n1814), .op(n1817) );
  nand2_1 U2070 ( .ip1(partialQ[3]), .ip2(n1815), .op(n1816) );
  nand2_1 U2071 ( .ip1(n1817), .ip2(n1816), .op(n1818) );
  nand2_1 U2072 ( .ip1(n1820), .ip2(n1819), .op(n1822) );
  nand2_1 U2073 ( .ip1(n1825), .ip2(partialQ[3]), .op(n1826) );
  nand2_1 U2074 ( .ip1(n1827), .ip2(n1826), .op(n454) );
  inv_1 U2075 ( .ip(n1898), .op(n1829) );
  nor2_1 U2076 ( .ip1(n1829), .ip2(n1828), .op(n1830) );
  not_ab_or_c_or_d U2077 ( .ip1(n1830), .ip2(n1899), .ip3(reset), .ip4(n441), 
        .op(n1831) );
  ab_or_c_or_d U2078 ( .ip1(n1833), .ip2(n588), .ip3(n1832), .ip4(n1831), .op(
        N317) );
  nand3_1 U2079 ( .ip1(n1850), .ip2(doB[3]), .ip3(n1854), .op(n1842) );
  mux2_1 U2080 ( .ip1(n1949), .ip2(n1835), .s(aAQ[7]), .op(n1948) );
  mux2_1 U2081 ( .ip1(n1920), .ip2(n1836), .s(aBQ[2]), .op(n1921) );
  mux2_1 U2082 ( .ip1(n1953), .ip2(n1837), .s(aBQ[7]), .op(n1904) );
  mux2_1 U2083 ( .ip1(n1929), .ip2(n1838), .s(aAQ[2]), .op(n1928) );
  ab_or_c_or_d U2084 ( .ip1(n1880), .ip2(doB[12]), .ip3(n1843), .ip4(n1839), 
        .op(n1840) );
  and2_1 U2085 ( .ip1(n1844), .ip2(doA[0]), .op(n1882) );
  mux2_2 U2086 ( .ip1(doA[6]), .ip2(doA[5]), .s(n1854), .op(n1887) );
  mux2_2 U2087 ( .ip1(doA[2]), .ip2(doA[1]), .s(n1854), .op(n1883) );
  nand2_1 U2088 ( .ip1(\mult/counterQ [2]), .ip2(doB[6]), .op(n1866) );
  nand2_1 U2089 ( .ip1(\mult/counterQ [2]), .ip2(doB[5]), .op(n1865) );
  inv_1 U2090 ( .ip(doA[6]), .op(n1884) );
  inv_1 U2091 ( .ip(doA[7]), .op(n1885) );
  inv_1 U2092 ( .ip(doA[2]), .op(n1878) );
  inv_1 U2093 ( .ip(doA[3]), .op(n1879) );
  inv_1 U2094 ( .ip(doA[4]), .op(n1876) );
  inv_1 U2095 ( .ip(doA[5]), .op(n1877) );
  inv_1 U2096 ( .ip(doA[1]), .op(n1875) );
  and2_2 U2097 ( .ip1(n1854), .ip2(doA[15]), .op(n1895) );
  nand2_1 U2098 ( .ip1(n1870), .ip2(doB[13]), .op(n1863) );
  nand2_1 U2099 ( .ip1(n1854), .ip2(doB[7]), .op(n1867) );
  nand2_1 U2100 ( .ip1(n1870), .ip2(doB[9]), .op(n1868) );
  nor2_1 U2101 ( .ip1(aBQ[4]), .ip2(n1945), .op(n1908) );
  nor2_1 U2102 ( .ip1(aAQ[4]), .ip2(n1945), .op(n1937) );
  nand3_1 U2103 ( .ip1(n622), .ip2(n1907), .ip3(aBQ[4]), .op(n1910) );
  nand3_1 U2104 ( .ip1(n622), .ip2(n1942), .ip3(aAQ[4]), .op(n1939) );
  and2_1 U2105 ( .ip1(n623), .ip2(aBQ[0]), .op(n1923) );
  and2_1 U2106 ( .ip1(n623), .ip2(aAQ[0]), .op(n1925) );
  and2_1 U2107 ( .ip1(aBQ[5]), .ip2(aBQ[4]), .op(n1901) );
  and2_1 U2108 ( .ip1(aAQ[5]), .ip2(aAQ[4]), .op(n1941) );
  nand3_1 U2109 ( .ip1(n1880), .ip2(\mult/counterQ [2]), .ip3(doA[0]), .op(
        n1881) );
  nand3_1 U2110 ( .ip1(n1880), .ip2(doB[0]), .ip3(n1892), .op(n1873) );
  nand3_1 U2111 ( .ip1(n1854), .ip2(n1851), .ip3(doB[15]), .op(n1864) );
  nand3_1 U2112 ( .ip1(n1854), .ip2(n1851), .ip3(doB[11]), .op(n1869) );
  nor2_2 U2113 ( .ip1(aAQ[4]), .ip2(aAQ[6]), .op(n1855) );
  nor2_2 U2114 ( .ip1(aBQ[6]), .ip2(n1945), .op(n1903) );
  mux2_1 U2115 ( .ip1(n1910), .ip2(n1909), .s(aBQ[5]), .op(n1911) );
  mux2_1 U2116 ( .ip1(n1913), .ip2(n1912), .s(aBQ[4]), .op(n4) );
  nor2_2 U2117 ( .ip1(aBQ[1]), .ip2(n1945), .op(n1916) );
  mux2_1 U2118 ( .ip1(n1919), .ip2(n1918), .s(aBQ[3]), .op(n5) );
  mux2_1 U2119 ( .ip1(n622), .ip2(n714), .s(aBQ[0]), .op(n8) );
  mux2_1 U2120 ( .ip1(n1925), .ip2(n1927), .s(aAQ[1]), .op(n9) );
  mux2_1 U2121 ( .ip1(n1932), .ip2(n1931), .s(aAQ[3]), .op(n11) );
  mux2_1 U2122 ( .ip1(n1935), .ip2(n1936), .s(aAQ[4]), .op(n12) );
  mux2_1 U2123 ( .ip1(n1939), .ip2(n1938), .s(aAQ[5]), .op(n1940) );
  mux2_1 U2124 ( .ip1(n1943), .ip2(n1946), .s(aAQ[6]), .op(n14) );
  nor2_2 U2125 ( .ip1(aAQ[6]), .ip2(n1945), .op(n1947) );
  mux2_1 U2126 ( .ip1(n1952), .ip2(n1951), .s(aAQ[8]), .op(n16) );
  mux2_1 U2127 ( .ip1(n1956), .ip2(n1955), .s(aBQ[8]), .op(n17) );
  mux2_1 U2128 ( .ip1(n623), .ip2(n714), .s(aAQ[0]), .op(n18) );
endmodule

